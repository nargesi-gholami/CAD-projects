module get_input(input clk, input [9:0] addr, input read_input, output reg [495:0] out);

reg[495:0] in[0:749];

assign in[0] = 496'b00010001_01110100_01101000_01100110_01101101_00000101_01101101_10110110_11111100_11111100_00000011_11111111_00011010_10110000_11111111_11111111_10111110_00111011_11111111_10111010_01000001_10101000_01001111_01111110_00110110_11111111_11100111_01101010_01111110_01111110_11000010_11111111_11001110_01011111_01001000_10100111_01001000_10011001_11111111_01011110_00001111_11110011_11111011_01000101_10010101_11111111_01001111_11111010_11010100_00111101_01100000_11101000_11111111_01111110_01101110_01111101_01011100_11011101_11111111_10011000_11110010_11111111;
assign in[1] = 496'b11111111_11111111_11111111_11111111_11111111_11101010_00001110_01110101_00111011_11001001_11111111_11111111_00110011_01111110_01111110_01111110_01001011_11111111_11110110_01110011_01111111_10000101_10111101_01111101_11011000_11111111_00111100_00001110_11111111_10011001_01111011_11100000_11111111_11111111_11111111_11111111_00110101_01000000_11111111_11111111_11111111_11111111_10111000_01111100_10100101_11111111_11111111_11111111_11110110_01011000_01101111_11111011_11111111_11111111_11111111_10110010_01111110_10110110_11111111_01011100_00111001_11111101;
assign in[2] = 496'b11111111_11111111_00001111_00101001_11111111_11111111_11111111_11111111_01001101_00101001_11111111_11111111_11111111_11111111_11110001_01111101_10001110_11111111_11111111_11111111_11111111_10001011_01100001_11110011_11111111_11111111_11111111_11111111_00110100_01010011_11111111_11111111_11111111_11111111_11100001_01110001_00010100_11111111_11111111_11111111_11111111_10000111_01111101_11100101_11111111_11111111_11111111_11111111_00101000_01111110_11111111_11111111_11111111_11111111_11111111_00101000_00110011_11111111_11111111_00101000_10110110_11111111;
assign in[3] = 496'b11111111_01011000_11101011_11111111_11111111_11111111_11111100_01100000_11101011_11111111_11111111_11111111_11111111_11101001_01011001_11111111_11111111_11111111_11111111_11111111_10011100_00101111_11111111_11111111_11111111_11111111_11111111_00101110_10110010_00000001_00100010_11100011_11111111_11000101_01111110_01101101_00100011_00110110_10011000_11111111_00000101_01101110_11100011_11111111_01000000_10011110_11101111_01101011_10111111_11111111_11111111_01010010_11100101_11111101_11010111_11111111_11111111_11011001_00001111_11111111_11111111_11111111;
assign in[4] = 496'b11100100_10111000_10100000_11100110_11111111_00010110_01110000_01111101_01111101_01101000_10110100_00111010_01111101_01000011_10010000_00010000_01111101_00111101_01111101_00111110_11111111_11111111_11111111_10001110_01101010_01110101_01111010_00111110_00011111_00011111_00101011_01100001_11101001_10010100_01000001_01000100_10010001_01010000_01000110_11111111_11111111_11111111_11111111_10111100_01111101_00001111_11111111_11111111_11111111_11111001_00111000_01101111_11000101_11111111_11111111_11111111_10110011_01111101_00110010_00110010_01111100_01000010;
assign in[5] = 496'b11011100_01001010_01010101_00101000_01101011_11110101_01011001_10000011_11111111_11110110_01011100_11111111_10100100_01011000_11111101_11111111_00100001_01010111_11111111_10011110_00101001_11101000_00100000_01011011_11010110_11111111_11001010_01111100_01110100_01001001_11101101_11111111_10000100_01100111_01001111_00001100_01010111_00010100_11101110_01110011_10010000_11111111_11111111_11111111_01001001_00001000_01110000_11001111_11111111_11111111_10011000_01101110_11010011_10100110_01101110_00111111_00101111_01100010_11001011_10010100_10010000_11100111;
assign in[6] = 496'b10110010_01111101_11001011_11111111_11111111_11111111_00111011_00100110_11111111_11111111_11111111_11111111_10101000_01111101_00111111_01001011_01001010_00001100_11011100_01110101_01111101_01000011_10000111_10000110_01011010_01000001_01101000_10100100_11111111_11111111_11111111_10111100_01111101_10100110_11111111_11111111_11111111_11111111_11001101_00100110_11111111_11111111_11111111_11111111_11111111_10101000_01011010_10010010_10111011_10111011_10111011_10001111_01110101_10101110_00101110_01111000_01011101_01001000_00111001_11111111_11111111_11111111;
assign in[7] = 496'b11111111_11001010_01101010_11110000_11111111_11111111_11111101_01000000_10000101_11111111_11111111_11111111_11111111_10111101_01100011_11110001_11111111_11110000_11111111_11111011_01001101_01000000_00011011_01001110_01111011_11111111_10101110_01110011_00100101_10101111_00101111_00101011_11111111_00111110_10010010_11111111_11010000_01101100_11100001_11000100_01101010_11110001_11111111_00110000_10011001_11111111_01001001_10101000_11111111_11000110_01011010_11110110_11111111_10000111_11111111_11111111_10000001_10000111_11111111_11111111_11111111_11111111;
assign in[8] = 496'b10011110_01001011_00011000_01000011_01100111_10101101_01011010_11010101_11111111_11000100_01111110_11101111_01110001_10101110_11111111_11111111_11110100_01110001_10110101_00101111_11111110_11111111_11111111_11111111_01011111_00110001_00000100_11111111_11111111_11111111_11101111_01110100_01100111_10000001_11111111_11111111_11111111_10100101_01100000_01100111_00000100_11111111_11111111_11011011_01101100_10010000_01000011_01100111_00001110_00101100_01110001_00101111_11111110_10100000_00110010_01111011_01111101_00101010_11110100_10111011_10101111_11111001;
assign in[9] = 496'b11111111_11111111_11111111_11111111_11110110_11111111_11111111_11111111_11101000_00011001_01100010_11111111_11111111_11111111_11011111_01010110_10001011_11110000_11111111_11111111_11111111_10000010_11000001_11100000_01000010_11111111_11111111_11111111_10011001_00011101_01100000_10011101_11111111_11111111_11111111_11011010_01101101_11001111_11111111_11101011_10101010_00010100_01100110_00000011_11111111_11111111_01001001_00001100_10110000_10111000_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111;
assign in[10] = 496'b11111111_11111111_11111111_11111111_11111111_11010000_10010001_11111111_11111111_11111111_11111111_10111111_00011011_11111011_11111111_11111111_11111111_11111111_00001001_11111011_11111111_11111111_11111111_11111111_10001010_11111111_11111111_11111111_11111111_11111111_11111111_00010111_11111110_11111111_11111111_11111111_11111111_11110111_10111000_10000010_00000111_10000011_10000100_00010111_00010101_00000010_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111;
assign in[11] = 496'b11111111_11111110_00111110_01111001_11000111_11111111_11111111_10010101_01111110_10001101_11111111_11111111_11111111_11100110_01100101_00101101_11111010_11111111_11111111_11111100_01001000_01010000_11111011_11100000_10011111_11111111_00000110_01111110_01010001_01011011_01111001_01111110_11000100_01111010_00101101_00010101_10001010_01101101_01000011_01001111_00011000_11111111_11111111_00011100_01101000_11011000_01010111_11111001_11111111_10101001_01110010_11001100_11111111_11001011_11111111_11111111_00110101_00000001_11111111_11111111_11111111_11111111;
assign in[12] = 496'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_11101110_10100110_00100100_00110111_11110111_10100001_00110001_01101101_01110111_01110111_01111010_01010010_01111100_00100101_11011000_11111111_11111111_11011011_01111010_10000111_11111111_11111111_11111111_11111111_10111110_01100100_11111110_11111111_11111111_11111111_10011100_01101010_01111101_00010011_11111111_11100111_00100100_01111101_10001100_01111010_01111101_00100001_01001101_01001100_11000101_11111111_00001100_01111010_01110100_00011111_11101100_11111111_11100111_11111111_11111111;
assign in[13] = 496'b11111111_11111111_11111111_11111100_11011111_11111111_11111111_10111010_00101001_01101000_01111110_11111111_11111111_11000000_01110001_00101011_00001011_11001101_11111111_11111111_00010011_10001111_11111111_11111111_11111111_11111111_11111011_01001111_11001001_11111110_10101101_11100100_11111111_11111111_10000011_00101000_00011011_01110010_11011111_11111111_11111111_11101010_01100111_01111000_10111000_11111111_10001011_00100011_01001100_01100101_11001111_11111111_11111111_01000000_01011110_01010011_11000001_11111111_11111111_11101100_11111111_11111111;
assign in[14] = 496'b11111111_11111111_10111001_10001001_11111000_11101111_10010111_01010011_01111100_01111100_00101010_11010010_01011100_01111100_01111101_01111100_01111100_01111100_01010010_01100010_10101110_00100001_01111010_00000111_01101100_01111100_10011100_00010111_01111011_10000011_00111111_00110111_01100110_01111101_01111010_00001110_00001011_01111011_10110100_11100000_10010101_11011110_10110100_01111100_10000100_11111111_11111111_11111111_11100110_01101111_00110101_11111001_11111111_11111111_11100101_01010101_01100001_11100110_11111111_01111100_00111011_11111111;
assign in[15] = 496'b11111111_11111111_11011000_01110101_00010011_11111111_11111111_11111111_00010000_01101100_11100100_11111111_11111111_11111111_10111101_01111001_10000110_11111111_11111111_11111111_11010100_01101101_00110011_11111111_11111111_11111111_11111100_01000111_01111101_01100001_01100000_00100100_11110010_01000101_01111100_01010010_00111101_01101111_01111101_00100100_01111100_10100001_11111111_11010110_01100110_00100100_01111010_10001011_11111111_11111111_01010100_01011101_11101011_00010110_11111100_11111111_11110101_01110100_10110011_11111111_11111111_11111111;
assign in[16] = 496'b00011011_01111101_01111101_01111101_01100100_00111100_01111101_00001011_11100011_10000010_01111101_00011001_01111100_10010000_11111111_11111111_11101100_01111101_01110011_00011111_11111100_11111111_11111111_11101100_01111101_01111101_11101010_11111111_11111111_11111111_10110101_01111101_01010111_11111001_11111111_11111111_11111100_01010010_01111101_01111101_11101011_11111111_11111111_10110010_01111101_01111101_01111010_10000010_11100100_11001000_01101010_01111101_01111010_00100110_01111010_01111101_01111101_01111101_01101000_10000001_10000001_10000100;
assign in[17] = 496'b11010001_10111101_11111111_11111111_11111111_11111111_10110111_00010100_11111111_11111111_11111111_11111111_11001100_00010100_01001001_10100100_11110110_11111111_11111111_10111000_00110111_01011000_01000011_10000110_11111111_11111111_11111111_11010010_00100011_10111010_00000100_11111111_11111111_11111111_11110111_00111110_11000011_00010101_11111111_11111111_11111111_11110010_01100101_11010000_11010100_11111111_11111111_11111111_11110101_01011010_11111111_11111111_11111111_11111111_11111111_11111111_01010010_11111110_11111111_11111111_01010101_11110111;
assign in[18] = 496'b11111111_11111111_11111111_11111111_11111111_00010101_11111111_11111111_11111111_11111111_11111111_11001011_01010011_11111111_11111111_10101011_00011100_01000000_11100101_01111101_00010010_01001001_01101110_00000110_01101011_11100101_01110100_00101011_10100011_11111001_11110000_01110000_11100101_00111110_11111111_11111111_11111111_10010110_01001110_11110000_10010111_11111111_11111111_11110111_01010000_10111011_11111111_11111111_11111111_11111111_10000111_01000101_11111010_11111111_11111111_11111111_11101100_01010111_11001100_11111111_10001100_00001111;
assign in[19] = 496'b01100010_01110001_01111101_01111101_01100001_01011010_10001000_11101111_11011111_10011000_00111011_10010100_01011000_11111111_11111111_11111111_11111111_11110100_00000111_00100100_11101100_11010111_10111100_11111111_11111111_10111001_01111101_01111101_01111101_01101100_11111001_11111111_10111101_01111000_00110111_10001010_11011010_11111111_11111111_01011011_00011000_11111111_11111111_11111111_11111111_11111111_01101111_10010000_11111111_11100110_10111100_00010110_01001001_10000110_01111000_01100011_01111000_01111101_01111100_10000001_10100011_10111100;
assign in[20] = 496'b11111111_10000101_00000000_11111111_11111111_11111111_11001101_01010101_11111010_11111111_11111111_11111111_11111111_00110011_10011110_11111111_11111111_11111111_11111111_11111111_01000110_10101111_11111111_11111111_11111111_11111111_11111111_00000000_01110111_01010101_11001101_11111111_11111111_11111111_11111101_00011011_01001110_11101101_11111111_11111111_11111111_00100000_01010000_11000101_11111111_11111111_11111111_11111111_00101000_01011110_01011101_00101101_11111111_11111111_11111111_11110101_10101111_10101111_11100000_11111111_11111111_11111111;
assign in[21] = 496'b11111111_11111111_11111111_11011011_01111010_11111111_11111111_11111111_11111111_00000001_01111011_11111111_11111111_11111111_11111111_10011011_01111110_00100011_11111111_11111111_11111111_10101011_01110011_01010111_11110111_11111111_11111111_11000111_01110011_01101011_11100111_11111111_11111111_11010110_01101010_01110011_11011000_11111111_11111111_11111100_01001000_01111110_10100100_11111111_11111111_11111111_10110100_01111110_00001101_11111111_11111111_11111111_11111111_01001000_01010001_11111111_11111111_11111111_11111111_11111111_11111111_11111111;
assign in[22] = 496'b11011101_11111111_11111111_11111111_11111111_00000000_01111011_11001110_11111111_11111111_11111111_11111111_11110101_01011110_10011101_11110010_10000110_01010100_11111111_11111111_00000110_01111001_01101100_01011000_10101101_11111111_10110011_01100011_01100111_01100000_00011110_01001010_10010001_01111101_10011111_11110011_10101010_10010111_11000011_01101110_10101100_11111111_11101001_11111110_11111111_11111111_01100001_10110011_00100110_01110101_10110101_11111111_11111111_01101110_01101100_00111110_10011011_11111111_11111111_11111111_11111111_11111111;
assign in[23] = 496'b11111111_11111111_00000100_01111100_10001110_11111111_11111001_00011001_01110111_10010001_11111110_11111111_11111111_00001000_01111001_10010010_11111111_11111111_11111111_11010011_01110111_00101010_11111111_11111111_11111111_11110010_01011100_01100100_11101110_11111111_11111111_11111111_10011000_01111100_10111110_11111111_11111111_11111111_11111111_01011101_00110101_11111001_11110111_10111101_00000010_00011101_01101001_01110011_01011101_01111101_01111011_01001110_10101110_10110100_10000001_10011101_11001011_11111111_11111111_11111111_11111111_11111111;
assign in[24] = 496'b11001000_01001011_01111110_01101011_00101100_00001010_01101000_10100101_11100100_10111000_00010100_11010100_01111101_10100101_11111111_11111111_11111111_11111111_10101110_01111110_11100100_11111111_11111111_11111111_11111111_11110100_01000110_01110010_01010010_01000101_00111000_11010111_11111111_11110111_10001100_01111110_00100110_00001101_11011110_11111111_11011000_01011111_10001001_11111010_11111111_11111111_11111111_00100110_00111001_11111111_11111111_11111111_11111111_11111111_10101000_01111011_00010011_10111000_11110100_10110100_00111001_01011111;
assign in[25] = 496'b11111111_11111111_11111111_11111111_11111111_10001111_11111111_11111111_11111111_11111111_11111111_00010000_10111110_11111111_11111111_11111111_11111111_11111111_01100001_11001001_11110010_11110010_11110010_11110010_10001110_01100001_01011100_01010011_01010011_01010011_01000000_01000111_01100001_11100100_11111111_11111111_11111111_11111111_01000010_01100111_11111111_11111111_11111111_11111111_11111100_01010000_01100010_11111111_11111111_11111111_11111111_11100100_01001000_00111001_11110100_11111111_11111111_11111111_11111100_11111111_11111111_11111111;
assign in[26] = 496'b10110011_01100001_01111101_01111101_10011001_11000000_01111101_00011110_10000101_01111000_11011110_11111111_10100100_01111101_10100000_00000010_01100000_11111111_11111111_11110001_01010000_01111101_01111101_10110000_11111111_11111111_11111111_11101100_01101100_01111101_01100110_11000101_11111111_11110010_01001000_00110011_11010001_01010100_01101111_11111010_01000100_01011111_11101101_11111111_11101101_01111101_00010001_01111101_10001101_11111011_10111000_01010000_01111001_01100101_01111101_01100001_01100111_01111101_01100000_10000001_10000001_11000100;
assign in[27] = 496'b10101011_01011011_01111000_01001101_01110110_10101111_01111010_00010101_11010011_11011011_00110011_11111111_00001101_01000000_11111001_11111111_11111011_11111011_11111111_00111000_00111010_11110101_11111111_11111111_11111111_11111111_10000011_01111101_01010101_10110001_11111111_11111111_11111111_11111010_10110001_01010001_01111011_00000011_11111111_11111111_11111111_11111111_11111111_10111110_01110011_11100101_00000010_11100011_11111111_11010000_00001110_01101000_10101111_01110110_01111000_01110101_01111001_00111111_11100101_10000010_10111100_11101100;
assign in[28] = 496'b11111111_10011010_01010000_11111111_11111111_11111111_11111111_00111101_10011101_11111111_11111111_11111111_11111111_11011100_01101000_11010100_10110000_11101100_11111111_11111111_10000001_00110001_01001110_00000000_01000111_11111111_11111101_01011010_01010110_11011111_11111111_01111010_11111111_10101010_01001111_11010110_11111111_11100101_01010011_11111111_00111000_11110001_11111111_11101011_01000001_10100010_11111111_01011111_11111110_11011101_01010111_10010110_11111111_11111111_00100101_01100100_01010011_10111100_11111111_11111111_11111111_11111111;
assign in[29] = 496'b11101000_00111100_01110000_00011010_00101001_11111111_10011001_01111001_11011100_11111111_11011101_11111111_11111111_10011001_01110011_11111100_11111111_10000111_11111111_11111111_11000110_01111011_00101010_00001111_01010010_11111111_11110011_10001101_01101101_01111101_00111001_11101110_10110100_01110010_01100100_10011000_00100000_01110010_11111111_01110001_01000111_11101011_11111111_10100100_01111110_11100110_01101011_11100110_11111111_11111000_00110110_01100110_11111111_01110101_10001100_10000010_01010100_01101100_10110110_10000010_10111000_11101110;
assign in[30] = 496'b11111111_11100011_01010000_01011101_11010000_11111111_11101110_01000111_01001000_11100001_11111111_11111111_11111001_00111101_01011111_11100010_11111111_11111111_11111111_00001011_01111101_10111110_11111111_11111111_11111111_11010101_01111101_00000100_11111111_11111111_11111111_11111111_00011111_01110010_11100101_11111111_11111111_11111111_11111111_01100000_00011101_11110100_11000111_10010101_00110111_01010111_01111000_01100101_01111000_01111100_01100001_10010001_11100010_10110101_10010100_10111010_11110010_11111100_11111111_11111111_11111111_11111111;
assign in[31] = 496'b11110010_10101110_10111010_11111011_11111111_11111111_11000000_10010010_01111000_01010011_00011111_11111111_11001010_00110000_01010010_01110111_10111001_01011000_11001010_01011100_10110010_11011110_01110110_11111000_01010000_01011101_11010010_11111010_00110100_10000110_11000110_01101110_01100101_11000011_01000000_00011001_11111111_00111011_10010011_10001111_00011011_10011000_11111110_10101010_00111110_11111011_11111111_11111111_11111111_11101101_01101100_11100001_11111111_11111111_11111111_11111111_00000010_00100101_11111111_11101101_01100110_11001110;
assign in[32] = 496'b11111111_11111111_11110101_01100001_10110100_11111111_11111111_11111111_10100010_01111110_11001001_11111111_11111111_11111111_11111000_01010111_01000111_11111111_11111111_10011111_11010011_00111101_01111101_00000110_11111111_11111111_11111111_11001010_01111100_00011110_11111110_11111111_11111111_11111111_00010100_01110011_11011110_11111111_11111111_11111111_11011010_01101001_00101111_11111111_11111111_11111111_11111111_10010000_01111100_11100010_11111111_11111111_11111111_11111111_01110011_00001100_11111111_11111111_11111111_11100011_11111111_11111111;
assign in[33] = 496'b11111111_11111111_10011011_01010100_11111111_11111111_11111111_11111111_10000101_01101111_11111111_11111111_11111111_11111111_11101111_01101100_01000110_11111111_11111111_11111111_10111010_01101111_01111101_00111110_11111111_11111111_11111111_11111010_01100011_01010111_11110100_11111111_11111111_11111111_10011111_01111101_10011001_11111111_11111111_11111111_11111111_01000011_01001011_11111111_11111111_11111111_11111111_11011101_01111101_10100101_11111111_11111111_11111111_11111111_10011110_01100111_11110010_11111111_11111111_10001001_11111111_11111111;
assign in[34] = 496'b11111111_11111111_11111111_11110101_10101100_00101011_11111000_11111111_10001111_01101100_01110100_10110111_01111110_11000110_00100001_01110100_00011010_11100111_10111110_01111001_01111100_01111101_00101011_10011111_00100011_11110010_01011010_01111100_01111101_01110110_01111000_00110000_10011101_01111000_10100010_10110110_10010101_11001010_11111111_01100101_00100011_11111111_11111111_11111111_11111111_11111111_01111101_11100000_11111111_10111110_10000111_11111111_11111111_00101001_11110100_00001010_01111101_00001101_11111111_01110011_10101111_11111110;
assign in[35] = 496'b11111111_11110100_00001001_01110100_01111100_11111111_11101010_01000010_01111101_01111110_01111011_11111111_11111111_11110101_01111100_01111100_01001110_10011111_11111111_11111111_11111111_01100111_01111100_11000110_11111111_11111111_11111001_00001100_01100001_01101011_10010101_11111111_11111001_00100101_01100001_11100001_00011000_00100100_11111111_00110001_01100001_11011101_11111111_10100001_01101001_11111111_01100001_11010111_11010110_10000011_01101101_10010011_11111111_01001011_01100110_01110000_00110011_10101101_11111111_11110100_11111111_11111111;
assign in[36] = 496'b00000010_01011000_01111100_01111100_00010101_00111010_00111000_10001001_10001001_00001011_01111100_01100000_00001010_11111011_11111111_11111111_11111110_00100101_00111101_11110111_11111111_11111111_11111111_11111111_10111110_00001110_11111111_11111111_11111111_11111111_11111111_00110000_00010110_11111111_11111111_11111111_11111111_11010011_01111100_01101011_11101101_11111111_11111111_11111111_00100110_01000110_00100011_00011101_11011010_11011111_10101011_01101111_11001001_11100110_00100100_01101010_01010001_01110110_10010000_00010010_01110111_00001001;
assign in[37] = 496'b11111111_11111111_11100100_01001101_01111001_11111111_11111111_11010000_01011100_01110001_10100101_11111111_11111111_11001111_01100101_01011101_11001111_11111111_11111111_11001000_01101111_01010000_11101000_11111111_11111111_11110100_01010101_01110000_11101011_11111111_11111111_11111111_00101010_01101010_11100101_11111111_11111111_11111111_11111111_01111100_10010011_11111111_11111111_11110001_11010000_10010010_01111100_01001110_00111101_01010100_01110110_01111001_00101001_10010001_10000001_10000010_10100010_10110110_11010110_11111111_11111111_11111111;
assign in[38] = 496'b01000100_01000000_11000101_11111111_11111111_01110100_01000101_00011111_01011001_11001111_11111111_11000111_00111100_11111111_11111111_11110010_01010000_11111011_00011011_10000111_11111111_11111111_10111110_01111110_11001101_10001011_01000010_10011001_00111110_01110010_00011010_10001110_11110101_01010001_01100101_00010100_11011011_10100100_00011011_11111111_11111111_11111111_11111111_11111111_00101011_00011011_11111111_11111111_11111111_11111111_10100100_01101000_11100000_11111111_11111111_10000011_00001011_01111010_00010110_00010011_01001101_10010010;
assign in[39] = 496'b11111111_11001011_01101100_01110000_11000011_11111111_11101011_01010101_01100101_11000101_11111111_11111111_11111111_00101001_01111100_11001101_11111111_11111111_11111111_11000000_01111101_00010001_10111011_11001111_11111111_11111000_01011101_01111101_01110111_01111101_01110101_10001111_10101001_01111101_00100101_11010000_11110100_00110100_00100101_01010000_01000111_11111111_11111111_11111011_01100000_10000100_10101110_00100110_11010111_11000001_00100001_01101110_11100101_11111101_00000010_01111110_01111110_00101101_11010111_11111111_11111111_11111111;
assign in[40] = 496'b11011110_11011100_01101100_01111100_10110010_11111111_11111011_10011001_01111101_00100000_11111111_11111111_11111111_11010001_01110110_00110101_11111000_11111111_11111111_11110011_01011001_01010001_11110111_11111111_11111111_11111111_00000101_01111010_10111001_11111111_11111111_11111111_11111010_01100010_01001111_11111111_11111111_11111010_11010010_11001111_01111110_10100111_11111110_11011000_10011000_01100110_10011101_01111101_00101100_01000010_01111101_01100001_00110011_10111001_01111110_01011110_00010010_10100010_11111100_11111111_11111111_11111111;
assign in[41] = 496'b00000110_01011000_00111011_00000001_11100011_10001111_01111011_10011110_11111011_11111111_11111111_11111111_00011111_01110100_11101001_11111111_11111111_11111111_11111111_11000011_01101111_01010011_11011000_11111111_11111111_11111111_11111111_11000101_01110001_01110000_10100100_11111111_11111111_11111111_11101110_00101011_01111100_00101011_11111111_11111111_11010101_01100100_01011010_10100110_11111010_11111111_11111111_00010110_01110010_11100010_11111111_11111011_11111111_11111111_11000011_01101100_01110001_01001101_01011010_11111101_10110010_10000010;
assign in[42] = 496'b11111111_11111111_11111111_00001010_01101111_11111111_11111111_11111111_11001011_01110110_00011101_11111111_11111111_11111111_11111101_01001110_01000100_11110111_11111111_11111111_11111111_10100101_01111011_11001001_11111111_11111111_11111111_11110000_01100000_00101010_11111111_11111111_11111111_11111111_10100000_01111101_11000110_11111111_11111111_11111111_11111110_01001001_00110111_11111101_11111111_11111111_11111111_10111000_01111100_10110011_11111111_11111111_11111111_11111111_00100010_00100111_11111111_11111111_11111111_10111101_11111111_11111111;
assign in[43] = 496'b11101110_00101110_01111100_01111101_01000100_11111100_00111100_01110111_00001111_00111111_01100111_11111111_00011011_01010101_11000110_11111111_00101110_01011111_11010110_01101111_11010110_11111111_11111111_00111100_01000001_00010011_01001111_11111111_11100101_11001000_01110111_10010001_00011010_10001000_11111111_00001111_01010011_01111100_11100011_00101100_10001000_10100110_01111101_01111101_10111010_11111111_00011010_01000000_01110110_01111101_01101000_11111111_11111111_10111011_01101011_01111101_01111101_00111001_11111111_10000010_11000101_11111111;
assign in[44] = 496'b11100111_11111111_11111111_11111111_11111111_01111101_11100111_11111111_11111111_11111111_11111111_11100111_01111101_11100111_11111111_11111111_11111111_11111111_11100111_01111101_11100111_11111111_11101010_10111010_11011010_11100111_01111101_00010000_00111110_00111111_00110010_01011010_11100111_01111101_00110100_11100100_11111111_11111111_11101100_11111110_00011110_00101010_11111111_11111111_11111111_10111111_11111111_11111111_00101010_00001110_10011011_00010011_01101111_11111111_11111111_11101111_10000001_10000001_10000001_11111111_11111111_11111111;
assign in[45] = 496'b01111100_01111101_01101011_00110011_11001010_01101001_01111100_01011110_01000011_01010101_01011011_11111111_01001001_01110010_11101110_11111111_11111111_11110110_11111111_11000001_01110111_00110011_00010010_11001011_11111111_11111111_11111111_11001101_01010000_01111101_01101010_11110010_11111111_11111111_11001101_01001111_01111100_00010110_11111111_11111111_10011011_01101100_01111101_00100001_11111000_11111111_11111111_01011011_01111100_00101001_11111001_11100111_11110000_11111111_11001000_01101100_01101000_01010100_01111010_11001101_00011011_01101011;
assign in[46] = 496'b11111111_11111111_11111111_10110000_11001101_11111111_11111111_11111111_11001010_01101000_11000010_11111111_11111111_11111111_11110001_01100101_10001111_11111111_11111111_11111111_11111111_00011011_00111011_10110010_00000011_00011010_00010110_00110111_01101011_00010100_01010011_01111100_11011001_11010110_01100000_00000000_00111100_01010011_10111110_11111111_00010110_01111110_01100000_00100000_11110100_11111111_11011000_01111110_01111110_10010010_11111101_11111111_11111111_11010100_00101011_11011011_11111111_11111111_11111111_11111111_11111111_11111111;
assign in[47] = 496'b11111111_11111111_11111111_11111111_11111111_10011011_11111111_11111111_11011000_00011000_01110011_10101111_01101001_11111111_10100101_01110011_01010101_10100100_11011000_01011111_01011111_01110011_10101111_11110110_00100010_10111001_01101001_01111101_01101001_01001011_01011111_00000100_01101001_00001110_11101100_10100101_10011011_11011000_11111111_00110111_11111111_11111111_11111111_11100010_11110110_11111111_00001111_11110110_10100101_00001110_01111101_11000011_11111111_01101001_01111101_01111101_01001011_10111001_11111111_11010111_11111111_11111111;
assign in[48] = 496'b11111111_11111111_11111111_11111111_11111111_10101111_11111111_11111111_11111100_10111100_01000000_10010100_01100000_11110110_10110001_01001110_01110101_00011011_11111111_01000001_01111101_01111101_01111101_00111011_00111111_11111111_01010101_01110110_00101101_00101101_00100111_11001000_10001101_01101111_10110000_11111111_11111111_11111111_11111111_01101001_10001011_11111111_11111111_11111111_11111111_11111111_01111101_11010101_10100010_10101111_00111000_11010000_11111111_01000100_01110100_01111001_01101011_00101100_11101100_10100110_11101100_11111111;
assign in[49] = 496'b11110011_00000010_01110101_01111100_01111100_11111111_00100000_01110101_10100000_10011010_01111100_11111111_11101000_01011101_00110000_10110010_01100100_00010011_11111111_11111101_01000011_01110010_01111010_10011111_11111111_11111111_11111111_10111001_01111110_01100110_11110110_11111111_11111111_11011111_01001101_01110010_01101111_00010110_11111010_10100101_01110100_01010111_11010001_01011111_01101011_11110000_01001100_01111100_01000110_00111010_01111011_01000100_11111100_01110011_00100010_00110100_00110100_10001000_11110000_11111111_11111111_11111111;
assign in[50] = 496'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111100_11111111_11111111_11111111_11111111_11111010_10110100_01010010_00100110_10110110_11111111_10101001_01010000_00111001_11111111_11010001_10000001_01101000_01111010_00010100_00110010_11111111_11111111_00000100_00001110_11011110_11001110_11111111_11111111_11111111_00111111_10110001_10000101_00101101_11010010_11111111_11111111_11001111_10001010_10110100_11100110_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111;
assign in[51] = 496'b01111110_11010101_11111111_11111111_11111111_11101000_01111111_11010010_11111111_11111111_11111111_11111111_11101000_01111110_11010010_11111111_11111111_11111111_11111111_11101000_01111110_11000000_11111111_11111111_11111111_01100011_01100110_01111110_01101110_01100011_01100011_01100011_10110101_10011110_01000001_01111110_10001101_10011110_10110101_11111111_11111111_11001001_01111001_00000100_11111101_11100001_11111111_11111111_11111111_00000001_01111110_01001000_01110110_11111111_11111111_11111111_11111001_10000010_00101111_11111111_11111111_11111111;
assign in[52] = 496'b01100111_01100101_10001100_11011101_11111111_01011011_10000111_10010000_01100000_01011010_11111111_11010010_01000100_11111001_11011000_10010101_01101110_11111111_11011100_00011000_11110010_01100101_00100100_01110100_11101100_11101111_01001011_00110011_00110111_00011100_01110011_11101111_11111111_11001111_11010110_11111111_00011111_01101110_11111111_11111111_11111111_11111111_11010010_01111000_00110010_11111111_11111111_11111111_11111111_10001011_01111100_10111011_11111111_11111111_11101011_10011100_01110111_00010001_11111111_01111110_01010111_11101001;
assign in[53] = 496'b11111111_11111111_10110111_00011000_11110100_11111111_11111111_10111100_01110110_01101100_11110100_11111111_11111111_11010110_01011111_10001011_11101110_11111111_10001100_11001001_01001101_01001001_11100111_11100111_10111010_00110111_01101100_01111101_01100111_01001011_01110001_01111101_11111111_10000111_01100111_11100111_10101111_01101100_00111111_11101111_01110110_00001100_00110100_01101100_10100100_11111110_10110100_01111110_01111000_00101111_11100100_11111111_11111111_11010000_01010110_00001010_11111110_11111111_11111111_11111111_11111111_11111111;
assign in[54] = 496'b10001110_01101010_01111101_01111101_01111101_00110001_01101111_00110011_10100001_11100011_10001111_01110111_01101111_11000001_11111111_11111111_11111111_11000000_01111101_10000011_11111111_11111111_11111111_11111111_11000000_01111101_10111101_11111111_11111111_11111111_11111111_00101101_01111101_10110110_11110110_11111111_11111111_10011100_01110110_01111101_01111101_01100111_11010011_00010000_01110100_01100011_01111101_01111101_01110110_01110001_01111101_01100101_11001010_01110011_01111101_01111001_01011001_00000101_11010111_11000110_11111111_11111111;
assign in[55] = 496'b11111111_11111111_00000001_10100110_11111111_11111111_11111111_11001111_01111001_11011010_11111111_11111111_11111111_11111111_00110100_00101011_11111111_11111111_11111111_11111111_11010011_01110111_10011111_10010010_00111001_01001010_01000011_01110100_01111110_01101001_01111110_01010111_10110011_10010001_01111101_00000010_01010111_00110000_11110101_11111111_10000110_01111101_01110110_00100011_11111111_11111111_11111010_01011011_01111110_00010011_11111011_11111111_11111111_11010011_01111110_00010100_11111100_11111111_11111111_11111010_11111111_11111111;
assign in[56] = 496'b00110110_01000100_01000101_00010011_11110101_01110101_01111101_01111101_01111101_01111101_00111101_00100111_01111101_00100001_10110010_00010000_01111101_01110100_01110100_01111101_11101001_11101000_11000001_01101000_10010101_00111001_01111101_00101010_01101100_01111101_01111101_01100111_10001101_01111101_01111101_01111101_01111101_01111101_01010111_11111001_01110000_01111101_01111101_01111101_00010111_11100010_11111111_01101101_01111101_01111101_01111101_10000100_11111111_11111111_00111000_01111101_01111101_01111101_10101000_01000110_01110111_10010111;
assign in[57] = 496'b11111111_11111111_10101010_01111000_10101111_11111111_11111111_11111011_01011111_00101000_11111111_11111111_11111111_11111111_00001001_01010110_11111011_11111111_11111111_11111111_10001100_01111101_10011010_11011101_11111111_11111111_11011000_01111000_01111101_01111101_01111000_10111001_11111111_00001001_01110011_10100101_11111011_00110001_10000001_10111001_01110011_11000011_11111111_11100111_01101001_10010110_00011101_00101000_11111111_11000011_01010000_01000001_11111011_10111110_01010101_01111101_01101110_10000001_11110001_11111111_11111111_11111111;
assign in[58] = 496'b11111111_11111111_11111111_11111111_11101101_11001100_11111111_11111111_11110011_00100110_01111100_01110000_00100010_11101000_00001111_01110110_01011100_10001100_00010100_01111110_01110110_01100101_10011101_11110110_10001011_11100101_01111010_01111110_01110101_00110101_01101010_01101111_10110001_01111110_10010111_10011000_00001000_00000001_11100001_01001000_00101000_11111110_11111111_11111111_11111111_11111111_01101100_10001111_11111111_11111111_11011010_00000100_11100010_00110001_01101000_00100001_00010101_01111001_01010000_01111110_00110000_10101000;
assign in[59] = 496'b11111111_00000111_01111110_00110111_11111111_11111111_11111111_01011011_01011001_01000000_11111111_11111111_11111111_11001011_01111110_01110001_10100111_11111111_11111111_11111111_10111100_01111101_00101010_11111111_11111111_11111111_11111111_00010010_01010101_00111011_11111111_11111111_11111111_10100010_00110111_11110110_00101101_10110101_11111111_11111111_00001110_10010101_11111111_10010110_00110111_11111111_11111111_00000001_10010001_11111111_10010010_01000000_11111111_11111111_11000000_01010101_10100011_01100011_10001011_10101100_10000001_11001110;
assign in[60] = 496'b11111111_11111111_11111111_10000011_01011110_11111111_11111111_11111111_11011000_01111010_00100000_11111111_11111111_11111111_11111101_00111100_01101110_11100011_11111111_11111111_11111111_10010100_01111100_10001000_11111111_11111111_11111111_10111001_01111010_00010000_11111110_11111111_11111111_11110100_01011000_01000110_11101011_11111111_11111111_11111111_00110000_01101010_11011101_11111111_11111111_11111111_11000111_01111100_10110000_11111111_11111111_11111111_11111111_01000100_00001110_11111111_11111111_11111111_11111111_11111111_11111111_11111111;
assign in[61] = 496'b11011010_00100100_01000001_11101000_11111111_11001100_01101011_00000110_11110110_11111111_11111111_11011101_01110001_10001111_11111111_11111111_11111111_11111111_11100101_01100010_00000011_11000110_11111111_11111111_11111111_11111111_11111100_10010011_01011101_00011001_11111111_11111111_11111111_11111111_11111111_00001001_00110101_11111111_11111111_11111111_11111111_11110101_01101101_11001100_11111111_11010111_11111111_11111111_11001001_01111011_11011010_11111111_10011000_11111111_11111111_11111111_00101011_00101010_00001010_11111111_11101010_10010000;
assign in[62] = 496'b11111111_11111111_01000101_01111101_10101100_11111111_11111111_11001000_01111101_01111101_00001101_11111111_11111111_11111111_00001101_01111101_01111101_11001000_11111111_11111111_11001000_01111101_01111101_00101001_11111111_11111111_11111111_10101100_01111101_01111101_10010000_11111111_11111111_11111111_01000101_01111101_01100001_11111111_11111111_11111111_11100100_01111101_01111101_00001101_11111111_11111111_11111111_10101100_01111101_01111101_11100100_11111111_11111111_11111111_10101100_01111101_01000101_11111111_11111111_01111101_10101100_11111111;
assign in[63] = 496'b10010000_00111010_01111100_01111100_01110101_01010100_01111100_01101000_00010011_00010011_00011001_01010100_01101100_10001010_11110100_11111111_11111111_11111111_01111100_10010001_11111111_11111111_11111010_11110011_11111111_01100001_01110111_00010000_00000110_01100001_01111101_11000011_11011010_01000010_01111100_01111101_01110001_00101011_11110010_11111111_00010100_01111100_00111010_11010011_11111111_11110010_11111111_01100001_01110110_11100000_11101101_10011101_01100100_11111111_00010001_01111100_01101000_01110010_01111100_00010111_01111110_01011110;
assign in[64] = 496'b11111111_11111100_00111011_10110110_11111111_11111111_11111111_10010101_01100110_11100011_11111111_11111111_11111000_11110001_01101100_10000100_11111111_11111111_11111111_00100101_01111100_01111110_01111100_01111010_01111010_11111111_11100100_01111011_10000110_11011001_01001001_01010101_11111111_11000110_01111110_11110100_11111111_01010110_10110110_11111111_00111100_00100000_11111111_11111111_10001000_11101110_11011111_01111000_11001110_11111111_11111111_11111111_11111111_10000100_01001111_11111111_11111111_11111111_11111111_11111111_11111111_11111111;
assign in[65] = 496'b00010011_11111111_11111111_11111111_11111111_00001011_10011011_11111111_11111111_11111111_11111111_11111111_00110111_10011011_11111111_11111111_11111111_11111111_11111111_00011111_10101110_11111001_10000110_01001000_01010110_11111111_00110011_00001011_01001010_00000111_11001101_11100010_11111111_01000010_01000110_10001001_11111111_11111111_11110000_11001110_01100010_00100011_11000101_11111111_11110100_00011110_01000001_00000110_01010000_10101110_01000000_00111101_10001111_10111001_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111;
assign in[66] = 496'b11111111_11111111_11111111_11111111_11111111_11111111_11001110_01011101_01111101_01111101_00010001_11111111_11011110_01101011_01111110_01111101_01111101_01111100_10101001_01101010_01011110_01111110_01111101_01110000_01111101_01101010_01100010_00011011_01111110_00011011_00011111_01111101_01111110_01111110_01101011_10000111_11110001_01011100_01110100_01111101_00110011_11100010_11111111_10010011_01111101_00011001_11110011_11111110_11111111_11111111_01010000_01111101_11001001_11111111_11111111_11111111_10110010_01111101_01000001_11111111_00010100_01101111;
assign in[67] = 496'b11011100_11111111_11111111_11111111_11111111_00110101_11011100_11111111_11111111_11111111_11111111_11111111_00110101_11000111_11110110_10110111_11010111_11111111_11111111_01001010_01111110_01111101_01111110_01110011_11001000_11111111_00110101_00000010_10110010_11000111_10010011_00010110_11111111_00111111_11011100_11111111_11111111_11111111_10011001_11111111_01111101_10011110_11111111_11111111_11111111_00010000_11010111_01111101_11000111_11111111_11111111_11111111_00010000_11010110_10110010_11111011_11111111_11111111_11111111_11111111_11111111_11111111;
assign in[68] = 496'b11111111_11111101_00101011_00110011_11100101_11111111_11111111_11001101_01111101_01111101_10111011_11111111_11111111_11111111_00011111_01111101_01111001_11100011_11111111_11111111_11010110_01111011_01111101_10000111_11111111_11111111_11111111_10011001_01111101_01110100_11100000_11111111_11111111_11110000_01010100_01111101_00010111_11111111_11111111_11111111_10111100_01111101_01110001_11001010_11111111_11111111_11111111_10111100_01111101_01001110_11111111_11111111_11111111_11111111_10111100_01111101_00001011_11111111_11111111_01111100_00001011_11111111;
assign in[69] = 496'b11111111_11111111_10011110_01101000_11111111_11111111_11111111_11111110_01010010_00000010_11111111_11111111_11111111_11111111_10011100_01111110_11000110_11111111_11000010_00000000_00111101_01110111_01111110_01001111_10100110_10010001_00000010_01001010_01111001_00001101_01100011_01011111_11111111_11111111_01100011_00110001_11111111_00110010_01001111_11111111_11000000_01111100_11000001_11110001_01110011_00010001_11111111_00010110_01101110_11111110_11111110_10100010_11110100_11111111_01001001_00100000_11111111_11111111_11111111_11011101_11111111_11111111;
assign in[70] = 496'b01101111_00010101_11111111_11111111_11111111_00101000_01000011_11111111_11111111_11111111_11111111_11111111_00101000_00011011_11111111_11111111_11111111_11111111_11111111_10110111_01101011_01100000_01001001_00001011_11100100_11111111_11111111_11100001_10000010_10000010_01010010_00001011_11111111_11111111_11111111_11111111_11111011_01010111_10101000_10010111_00001100_10011011_11101101_10111000_01101110_11101010_11001010_00001001_01010011_01010010_01011001_00010010_11111111_11111111_11111111_11111000_01100101_01011101_11100010_11111111_10111000_10111111;
assign in[71] = 496'b10010010_01011111_01111110_01001001_00001001_11001010_01111110_01100101_00100101_00110110_01110111_11111111_00010010_01111010_11011100_11111111_11111111_11011110_11111111_00110000_01110110_11100010_11111111_11111111_11111111_11111111_11010000_01110110_01110000_01011000_00101011_10001110_11111111_11111111_11010000_00101111_01111110_01111110_01111110_11111111_11111111_11111111_11111111_11110011_01010010_01010101_11100000_10101000_10000100_00101101_01110000_01111101_10001101_01111110_01111110_01111110_01111110_01101000_00001010_11110111_11110111_11111011;
assign in[72] = 496'b11111111_11111111_11111111_00100001_10010001_11111111_11111111_11111111_10111100_01010100_11111000_11111111_11111111_11111111_11101100_01100110_10010101_11111111_11111111_11111111_11111111_00001111_01100000_11101110_11111111_11111111_11111111_11101010_01101101_00000000_11111111_11111111_11111111_11111111_10100111_01111101_11100100_11111111_11111111_11111111_11111111_00111110_01100111_11111111_11111111_11111111_11111111_11111101_01100010_10001011_11111111_11111111_11111111_11111111_10101110_01110011_11010111_11111111_11111111_10110010_11111111_11111111;
assign in[73] = 496'b10011001_01101000_00011011_00111001_11100000_11101001_01110010_11010001_11111111_00000000_10101100_11111111_10101100_01001110_11111111_11111111_11110010_11110010_11111111_10101100_01000101_11111111_11111111_11111111_11111111_11111111_11000010_01110100_10111101_11010110_10110101_11111111_11111111_11111111_10001110_01001110_01111101_00010110_11111111_11111111_11111111_11111111_00101110_00100011_11111111_11111111_11111111_11111111_10010010_01001101_11110101_11111111_11111111_11111111_11111111_00001010_01101000_00011010_00110011_11111101_10100111_10000001;
assign in[74] = 496'b11111111_00101110_01111110_01111110_01110110_11111111_11001111_01111011_01001011_01111110_01110111_11111111_11111111_11011111_01111111_01111011_01101010_10110001_11111111_11111111_11101100_01110001_01111110_10001111_11111111_11111111_11100111_01001101_01100110_01111101_00101111_11111011_11011011_01010110_00110101_11110010_10010101_01111110_10011001_01000011_01111001_11100110_11111110_10001011_01111110_00001001_01100010_01111110_00000001_01000110_01111110_01011010_11011111_10100111_01111110_01111001_01000010_10101000_11110100_11101101_11111111_11111111;
assign in[75] = 496'b11111111_11111111_11110100_01011001_00101110_11111111_11111111_11111111_11001001_01111101_00111111_11111111_11111111_11111111_11111011_00111010_01111101_10000101_11111111_11111111_11111111_00011001_01111101_01000001_11111101_11111111_11111111_11001101_01110100_01111101_10010001_11111111_11111111_11111111_10101011_01111101_01100111_11101001_11111111_11111111_11110001_01100110_01111101_10111010_11111111_11111111_11111111_10101011_01111101_00111011_11111010_11111111_11111111_11111111_01010010_01101010_11100110_11111111_11111111_00100111_11110011_11110100;
assign in[76] = 496'b11000000_00101110_10010111_11111111_11111111_11111111_11111000_11000001_10010100_11111111_11111111_11111111_11111111_11111111_10000110_00011111_11000001_11111111_11111111_11111111_11111010_01000111_00111010_01000011_11010101_11111111_11111011_00101101_01000110_11111111_10000010_11001000_11111011_00011001_00111101_10011010_11111111_00100010_11101000_11100111_11101000_00111001_11110101_11111111_00100100_11101000_11111111_10111001_00000110_11111111_11111111_00100100_11101000_11101111_10000110_11110101_11111111_11101100_01011110_11111111_11111111_11111111;
assign in[77] = 496'b00101101_01110000_00100111_11001101_11111111_11001101_01111101_00011011_01010010_01111000_11110001_11111111_11111111_00111010_01011100_00001000_01111110_11010110_11111111_11111111_11100100_01010110_01111110_01100001_11111111_11111111_11111111_11011111_00111110_01111110_01110110_10101011_10001100_00101101_01111011_01011010_10001101_00111110_01111101_01111101_00101000_10100011_11110000_11111111_11111111_00110011_00110010_10100000_11010010_11010110_10111110_10001001_01100010_10000001_00110111_01110001_00111001_00110010_10000001_11111111_11111111_11111111;
assign in[78] = 496'b11101001_01100111_01110100_11010001_11111111_11111111_11110010_01010100_01001111_10011100_11111111_11111111_11111111_11111111_00110111_01111110_10100100_11111111_11111111_11111111_11111111_10110100_01111110_10101111_11111111_11111111_11111111_11101100_01100011_01110110_10011000_11111111_11111111_11111100_00110011_00100010_10001101_00111111_11111110_11111111_10001001_00111101_11111110_10011011_01111110_11110100_11100111_01110001_00110001_00111001_01110000_10000111_11111111_00110101_01100110_00110101_10100010_11010100_11111111_11001110_11111111_11111111;
assign in[79] = 496'b11111111_11111111_10100001_01110110_11101001_11111111_11111111_11111111_01000001_01110100_11101100_11111111_11111111_11111111_11101010_01111101_01001001_11111111_11111111_11111111_11111111_00011001_01111101_10011111_11111111_11111111_11111111_11110011_01101001_01100011_11110100_11111111_11111111_11111111_10011001_01111110_10000010_11111111_11111111_11111111_11110010_01100110_01110100_11110110_11111111_11111111_11111111_10111111_01111101_10001111_11111111_11111111_11111111_11111111_00011010_01011010_11111000_11111111_11111111_00000000_11111111_11111111;
assign in[80] = 496'b11101101_00000010_01111001_01111101_01111101_11011100_01100001_01111101_01000101_10011010_01111101_11101011_01010100_01100101_11000100_11111100_11010101_01111101_00011001_01100101_11011010_11111111_11111111_01000101_01101111_01101010_10111000_11111111_11111111_11010101_01111100_10000010_01010010_11111111_11111111_11111111_00101000_01110100_11101101_01010010_11111111_11111111_00000010_01111101_00000101_11111111_01110110_10111010_10110110_01110111_01111101_11110011_11111111_01010101_01111101_01111101_01111101_00110100_11111111_10000001_10111100_11111101;
assign in[81] = 496'b11110110_00001010_01001001_10000100_11101011_11111111_00010110_01111001_00111101_01010100_01111101_11111111_11110001_01110110_00010101_11111111_11111111_11011001_11111111_11111111_01011010_00111111_11101111_11111111_11111111_11111111_11111111_11000000_01111000_01010111_00110100_00011001_11111111_11111111_11111111_10011111_01100011_01111101_01110010_11111111_11111111_11000011_11001011_00010011_01111101_00100111_00110100_01111100_01111100_01111101_01111100_01001011_11101010_01001000_10000001_11010000_11110101_10110001_11100110_11111111_11111111_11111111;
assign in[82] = 496'b11111111_10010000_00001100_11111111_11111111_11111111_11111111_10011001_00101110_11111111_11111111_11111111_11111111_11111111_00001101_00010000_11111111_11111111_11111111_11111111_11111111_00010110_10000001_11111111_11111111_11111111_11111111_11111111_00110011_10110000_11111111_11111111_11111111_11111111_11111111_01011101_11011001_11111111_11111111_11111111_11111111_11100100_01111000_11100111_11111111_11111111_11111111_11111111_11100100_01110000_11111111_11111111_11111111_11111111_11111111_11100100_01101011_11111111_11111111_10110000_00101111_11111111;
assign in[83] = 496'b11111111_11010001_01101111_01101111_11110000_11111111_11111111_01010000_01111111_00010000_11111111_11111111_11111111_11000000_01111111_01010000_11111111_11111111_11111111_11111111_01010000_01111111_01000000_01101111_01111111_11111111_00100000_01111111_01111111_01011111_00010000_01111111_00000000_01111111_01101111_10110000_11111111_10110000_01111111_01111111_01111111_11110000_11100000_10100000_01101111_01010000_01100000_01111111_01000000_01101111_01111111_00000000_11110000_00000000_01111111_01000000_00100000_11000000_11111111_11111111_11111111_11111111;
assign in[84] = 496'b11111111_11111111_00000100_01110010_11110111_11111111_11111111_11111111_10000001_01111100_11110100_11111111_11111111_11111111_11110001_01111010_00110010_11111111_11111111_11111111_11111111_00001011_01110100_11010011_11111111_11111111_11111111_11110001_01101100_00111111_11111111_11111111_11111111_11111111_10100101_01111101_10011111_11111111_11111111_11111111_11111111_00100100_01111101_11101011_11111111_11111111_11111111_11111011_01100110_01110000_11111111_11111111_11111111_11111111_11111110_01010111_01100000_11111111_11111111_01001100_10011101_11111111;
assign in[85] = 496'b11111111_11111111_11111111_11101000_10100011_00110100_00001010_10111001_10000100_01110011_01111100_11100100_10101000_00000111_01111011_01001111_10000011_11001010_11111111_11111111_11001110_01101101_11100111_11111111_11111111_11111111_11111111_00100000_10000100_11111111_11111111_11111111_11111111_11111111_01110001_11011110_11111111_11111111_11111111_11111111_11111111_01111100_11110000_11111111_00011100_10111111_11111111_11111111_01101110_11101011_11111111_00100111_10110001_11111111_11111111_00011001_10000110_11110001_01100100_10110001_01100011_01001101;
assign in[86] = 496'b10011010_01100110_01111101_01111101_01111101_10101100_01111010_00111100_10101111_11111000_10000001_00001101_01111101_00000011_11111111_11111111_11111111_10111110_01110110_01010111_11111101_11111111_11111111_11111111_00010110_01111101_00000111_11111111_11111111_11111111_11011000_01111010_01111101_10001010_11101010_11101001_10001010_01111001_01111001_01111101_01110010_01101111_01110000_01111101_01111100_10000010_01111101_01111101_01111101_01111101_01111101_10000010_11111111_00011011_01001110_01111010_01111001_10000010_11111111_10011100_10101011_11111111;
assign in[87] = 496'b11111111_11000111_01101110_11110000_11111111_11111111_11111111_00111011_00001100_11111111_11111111_11111111_11111111_11000110_01111101_11100111_11111111_11111111_11111111_11111100_01001111_00100000_11100111_10111011_00000000_00110101_01001010_01111110_01110000_01111110_01111110_01011011_10100100_01111110_10001101_11100010_00001000_01110001_11100001_00110110_00110100_11111111_11111111_00011101_01000010_11101011_01111110_11011100_11111111_11111111_10110000_01101000_10110011_00101010_11111111_11111111_11111111_11111111_11111101_11111111_11111111_11111111;
assign in[88] = 496'b11111111_11111111_10011000_00011000_11111111_11111111_11111111_11101110_01100001_10111010_11111111_11111111_11111111_11111111_00011001_01000011_11111110_11001011_11111111_11101101_00000000_01111100_00111010_01100001_01111110_00010011_01111001_01111110_01010100_01011001_01111110_01010111_11101011_01101010_00111010_11110000_01011111_01011000_11100110_10001001_01110010_11001110_10111000_01111010_11011101_11111111_01111001_10010110_11111111_10101111_01011011_11111111_11111111_00111011_11110110_11111111_11111001_11110101_11111111_11111111_11111111_11111111;
assign in[89] = 496'b11111111_11111111_10111011_10000010_10000010_11011010_00010000_01001100_01001101_00110000_01000111_00101011_01001110_10011111_11101010_11111111_00100010_11000101_01111000_00001001_10011010_10011001_00110101_01101010_10011010_00010100_01000111_01000111_00111001_10010101_10110000_01101110_11111111_11111111_11111111_11111111_10101010_01110000_01100100_11111111_11111111_11111101_10001001_01111101_01010110_11100011_11111111_11100101_01000001_01111110_00101100_11111000_11111111_10111100_01101001_01110110_10000010_11111111_11111111_11001001_11111111_11111111;
assign in[90] = 496'b11111111_11111111_11000000_01111001_10011010_11111111_11111111_11100100_01011101_01001110_11111101_11111111_11111111_11110101_01001110_01101010_11101011_11111111_11111111_11111111_00100101_01111001_10111001_11111111_11111111_11111111_10110101_01111101_00000011_11111111_11111111_11111111_11101011_01100011_01011110_11111111_11111111_11111111_11111111_00110001_01110001_11000001_11100000_10111010_00010011_00111011_01111001_01111101_01110111_01101100_01001100_01101111_01100110_10001011_10011011_11101000_11111010_11111111_11000000_11111111_11111111_11111111;
assign in[91] = 496'b11111001_01001000_01110010_11010101_11111111_11111111_10011011_01111101_10000010_11111111_11111111_11111111_11010101_01110111_01001111_11110100_11111111_11111111_11111111_00110100_01100110_11101010_11111111_11111111_11111111_11000100_01111000_00000000_11111111_11111111_11111111_11101111_00010011_01110110_11100010_11111111_11111111_11101101_01000110_01111010_01010000_11111111_11100000_00000011_01101110_01111101_01111101_01111010_01110100_01111010_01111101_01111101_00111101_10101011_10000001_10000001_10011000_11100110_11100011_11111111_11111111_11111111;
assign in[92] = 496'b11111111_11111111_11011101_01100011_00011110_11111111_11111111_11111111_00011000_01111110_10100100_11111111_11111111_11111111_11001001_01111110_00110101_11111101_11111111_11111111_11111110_01010010_01110010_11010110_11111111_11111111_11111111_10011100_01111110_00011101_11111111_11111111_11111111_11111001_01001101_01101011_11101101_11111111_11111111_11111111_10111010_01111110_00011101_11111111_11111111_11111111_11111111_00111001_01111110_11000111_11111111_11111111_11111111_11111111_00110000_01010001_11110101_11111111_11111111_00001010_11111111_11111111;
assign in[93] = 496'b11111111_11111111_10100010_01111100_10101010_11111111_11111111_11011101_01110100_00110011_11111111_11111111_11111111_11101001_01100010_01001101_11110100_11111111_11111111_11111111_00111011_01110100_11011111_11111111_11111111_11111111_00000000_01110100_11000000_11111111_11111111_11111111_10100111_01111100_10001111_11111111_11111111_11111111_11111111_01100111_00101110_11111110_11111111_11111111_11101110_11111111_01111101_01110010_01010110_01100001_01101011_01110101_01100011_10000001_10000001_10001100_11001010_11001011_10011000_11111111_11111111_11111111;
assign in[94] = 496'b01011010_01001100_01011111_10111110_11111111_10011010_01011010_11111011_01000001_10111110_11111111_11111111_11001101_01110011_00010011_01001011_11111011_11111111_11111111_11111111_10010101_01111101_01001011_11011000_11111111_11111111_11111011_00011000_10001011_00001001_01101110_00110001_11111111_10000001_00100011_11111111_11111111_11110001_00110110_11101100_01110011_11011101_11111111_11111111_11000100_01010101_10000111_00100111_11110110_00100010_01100100_01100000_10011111_10100101_01010101_10000010_01010000_01111101_10101010_10000001_10101010_11001000;
assign in[95] = 496'b11111111_00011101_01111010_01110011_01101000_11111111_11101101_01110110_10011010_11111111_01111101_11111111_11111111_11100001_01111101_11100000_10010000_00111111_11111111_11111111_11111000_01100111_01010010_01011000_11011001_11111111_11111111_11101110_01011111_01111000_11001100_11111111_11111111_11001000_01100001_01110111_01110111_11101101_11111111_11010100_01110100_01001001_11000101_01111101_11001011_11111111_01110100_00111101_11101110_00011110_01010100_11111111_11111111_00110000_01111001_01110011_01110100_10011011_11111111_10010011_11100010_11111111;
assign in[96] = 496'b11111111_11111111_11111111_01011110_00101011_11111111_11111111_11111111_10101001_01101000_11011110_11111111_11111111_11111111_11010011_01100010_00101101_11111001_11111111_11111111_11111110_00011001_01111001_11100001_11111111_11111111_11111111_11000010_01111110_00000110_11111111_11111111_11111111_11111001_01001010_01101011_11011010_11111111_11111111_11111111_10111100_01111001_00101110_11111111_11111111_11111111_11111111_00111001_01111001_11000111_11111111_11111111_11111111_11111111_01000010_01001101_11110110_11111111_11111111_11001101_11111111_11111111;
assign in[97] = 496'b11111111_10110011_10000110_11100111_11111111_11111111_10100011_00101010_10011000_00101100_11111111_11111111_11111111_01011100_11100011_11001111_00101010_11111111_10101101_00111011_01110101_00000001_01010101_10111010_11111111_11111111_11011010_01100000_10000011_11001110_11111111_11111111_11111111_11111111_00001000_10101101_11111111_11111111_11111111_11111111_11111111_11001110_01000110_11111111_11111111_11111111_11111111_11111111_11111111_00010111_10101001_11111111_11111111_11111111_11111111_11111111_11101100_01001111_11100101_11111111_11111111_10111001;
assign in[98] = 496'b01110001_01101101_00010111_10000110_00010000_01111101_00110011_11100001_11111111_11111111_11111111_00101001_01111101_11001110_11111111_11111111_11111111_11111111_10101011_01111101_10101000_11111111_11111111_10111111_00101111_11111111_00101100_01110011_01001110_01001110_01111100_01111101_11111111_11111111_10111010_00011000_00101001_10001010_01111101_11111111_11111111_11111111_11111111_11111111_11001000_01111101_11100101_10100110_10000111_10000111_00011001_01100000_01111101_01111110_01111110_01111110_01111110_01111110_01111110_11111111_11111111_11111111;
assign in[99] = 496'b11111111_11111111_11010100_01110010_10011101_11111111_11111111_11111111_00100000_01111100_11001100_11111111_11111111_11111111_11011111_01111010_01001101_11111111_11111111_11111111_11111111_00000110_01111101_10100011_11111111_11111111_11111111_11111011_01100010_01001111_11110001_11111111_11111111_11111111_10011110_01111100_10000111_11111111_11111111_11111111_11111111_01000110_01110100_11100010_11111111_11111111_11111111_11001001_01111101_00100011_11111111_11111111_11111111_11111111_10111111_01111100_11010011_11111111_11111111_01011011_11111101_11111111;
assign in[100] = 496'b01001101_11111111_11111111_11111111_11111111_11100010_01010100_11111111_11111111_11111111_11111111_11111111_11100010_01010100_11111111_11111111_11111111_11111111_11111111_11100010_01010100_11111010_10010001_01010000_00110111_11111111_11001011_01010100_01001000_00001010_11110010_10100111_11111111_10011111_01110111_10101100_11111111_11111111_00000010_11111111_10011101_00110110_11111111_11111111_10101100_01010001_11111111_00000111_10000111_11110100_00000010_01000010_11100110_11111111_11010110_01000100_01100000_00000100_11111110_11111111_11111111_11111111;
assign in[101] = 496'b11100001_01000001_01110101_01101011_01110000_10001100_01010111_10001100_11011001_11111111_11110001_10110011_01111010_10101010_11111111_11111111_11111111_10111001_01101011_00100000_11111111_11111111_11111111_11101111_01011011_01111101_11100001_11111111_11110100_10110001_00101111_01111100_01111110_11111111_11111111_00110100_01111110_01111101_01001010_01111101_10110011_10111000_01100010_01111101_01100001_11101110_01111101_01110101_01100101_01111100_01111101_10101000_11111111_01000111_01111100_01111101_01111100_01110011_11100110_10000001_10100001_11101001;
assign in[102] = 496'b10111110_10000001_10000010_10010100_11110001_01000100_00111100_00010101_00100000_01100111_01011110_01101110_11010111_11111111_11100101_10010001_11100101_01101111_01111011_00011000_10001101_00110011_01101100_11010111_01101111_00100111_01111101_01101111_00111100_10101111_00000111_01110010_11111110_11101111_11110110_11111111_11001010_01111001_00101110_11111111_11111111_11111111_11010101_01100111_01100010_11101101_11111111_11111111_11000010_01101000_01100010_11010101_11111111_11111111_11000111_01111000_01001101_11101101_11111111_01010111_11100100_11111111;
assign in[103] = 496'b10011110_11111111_11111111_11111111_11111111_00010100_10011110_11111111_11111111_11111111_11111111_11111111_00010100_10010100_11001100_10111110_11110111_11111111_11111111_00000000_01110111_10001110_10000001_01000100_11011010_11111111_00000000_00101101_11111111_11111111_11001000_00111110_11111111_00010001_10001000_11111111_11111111_11111110_01100001_11111111_10011010_00010000_11111111_11111111_11111010_01101101_11111111_11101110_01011001_11000001_11011100_00100101_00101110_11111111_11111111_10111100_00111111_01100111_00010110_11111111_11111111_11111111;
assign in[104] = 496'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_00111000_00111000_00100001_00111000_00111000_00111000_00111000_00110000_01100110_01111110_01111010_00101110_10001001_01110100_11111111_00011110_01100111_11101010_11111111_11100011_01111110_11100001_01111100_00000011_11111111_11111111_11100011_01111110_00000011_01111110_11101101_11111111_11111111_11111101_01000110_01011001_01000111_11111110_11111111_11111111_11111111_11111111_01111110_10100111_11111111_11111111_11111111_11111111_11111111_11111111_11111111;
assign in[105] = 496'b11111111_11111111_11111111_10010001_00100001_11111111_11111111_11111111_11011011_01110011_10110111_11111111_11111111_11111111_11111111_01001110_00111001_11111111_00000111_10101111_11111000_10101001_01111000_11011010_11111111_11111000_10011010_01001111_01100101_00000011_11111111_11111111_11111111_11111111_00010110_01010011_00100000_11010110_11111111_11111111_10101100_01111000_11001100_11111111_11111111_11111111_11111111_10110011_01011101_01010000_01100010_00111010_00110010_11111111_11111111_11111100_11011111_11000011_11000001_11111111_11111111_11111111;
assign in[106] = 496'b11111111_11111111_11100111_11010000_00000001_11111111_11000110_01000000_01111000_01011111_00100001_11101110_00011010_01111110_01000001_11001111_11111111_11111111_00110110_01110000_10011101_11111111_11111111_11111111_11111111_01111110_10101011_11111111_11111111_11111111_11111111_11111111_01111110_10000010_11001010_10101001_00001001_00101010_01010010_10001010_01110010_01111110_01110110_00101110_10101101_11101101_11111111_00101001_01111110_01111011_00110100_10010100_11111111_11111111_11110010_10011000_10000101_00101111_00011101_11111111_11111111_11111111;
assign in[107] = 496'b11111111_11111111_11010001_01010010_01000011_11111111_11111111_11111111_00101010_01111101_10010000_11111111_11111111_11111111_11111111_00110110_01100101_11101100_11111111_11111111_11111111_10110001_01111101_10010101_11111111_11111111_11111111_11111001_01010110_00111100_11111111_11111111_11111111_11111111_10001001_01111100_11010001_11111111_11111111_11111111_11010111_01101111_00001010_11111111_11111111_11111111_11111111_00101010_01011101_11111000_11111111_11111111_11111111_11101111_01110000_00110110_11111111_11111111_11111111_00011111_11111111_11111111;
assign in[108] = 496'b11111111_11100100_11010001_11010001_11101011_11111111_11010110_01101000_01111110_01111110_01111100_11111111_11111111_00100000_01101101_10100000_10101111_00010110_11111111_11010011_01111100_10111010_11111111_11111111_11111111_11111111_11010100_01111110_10110100_11111111_11100101_11001101_11111111_11111110_00011010_01101111_01100100_01111001_00111011_11111111_11111111_11111111_00011000_01111110_00111011_11011010_11110110_11101010_10100001_01010100_01111110_11011011_11111111_01111010_01111010_01100100_01000110_00001011_11111111_11111111_11111111_11111111;
assign in[109] = 496'b11111111_11100010_00100111_01010101_10000001_11111011_00011101_00111100_10100101_11111011_11111111_11111111_00100010_10001011_11111011_11111111_11111111_11111111_11111111_00101101_11111111_11111111_11111111_11111111_11111111_11111111_11000100_00100010_11100010_11111111_11111111_11111111_11111111_11111111_11011101_10000111_00001001_10111001_11110001_11111111_11111111_11111111_11111111_11110001_00100111_01100100_11111111_11100111_10111110_00000100_01010101_00011001_11010111_00110001_00111011_00100010_10011011_11110001_11111111_11111111_11111111_11111111;
assign in[110] = 496'b10100110_01111000_00100101_01101110_10110011_11111111_00101100_00110000_11111111_10000001_01001111_11111111_11111111_00101100_00011111_11111111_10010010_00110011_11111111_11111111_00001101_01110011_11011011_01010100_10101010_11111111_11111111_11101101_01101001_01110001_00101000_11111110_11111111_11111111_11111111_01011100_01111110_11101100_11111111_11111111_11111111_00101000_01101110_01110011_10100110_11111111_11110110_00010100_01101100_11011110_00010010_00111110_11111111_01010110_00011111_01001000_01100010_01100010_01010011_11111111_11101101_11000101;
assign in[111] = 496'b11111111_11111111_11111111_10100011_11111111_00001011_00010101_10111010_11010010_01000101_11111111_11101001_11100100_11110011_00101100_01010000_10001001_11111111_11111111_11111111_11111111_10111100_01101111_11010001_11111111_11111111_11111111_11111111_11111110_00101010_11111111_11111111_11111111_11111111_11111111_11000011_10001111_11111111_11111111_11111111_11111111_11111111_00010101_11010010_11111111_11111111_11111111_11111111_11111111_00111110_11111111_11111111_11111111_11111111_11111111_11100110_00101010_11111111_11111111_11100001_00001111_11000100;
assign in[112] = 496'b11110110_00000001_01011010_01010011_11010111_11111110_00101000_01111110_01101100_01100101_01101011_11111111_10011101_01111101_00010000_11111111_10111111_01111101_11111000_01011100_00101111_11111111_11111111_00110000_01111101_10111110_01111110_10000110_11111111_10111010_01110110_00111101_10111111_01111101_10001110_11111111_00101001_01111010_11001011_11000001_01111101_10010111_11010111_01111101_00110010_11111111_11111110_01011001_01000001_00011111_01111101_10111111_11111111_11111111_01001101_01111101_01111110_00111111_11110110_01010011_01000011_11100110;
assign in[113] = 496'b00110010_11111111_11111111_11111111_11111111_10110101_00110010_11111111_11111111_11111111_11111111_11111111_10110101_00110010_11111111_11111111_11111111_11111111_11111111_10111010_00110010_11111001_10100000_00011000_00001001_11111111_11100111_01100111_01010000_00101000_10000001_00010011_11111111_10011011_01011101_11100100_11111111_11111111_11111111_11101010_01110001_00100011_11111111_11111111_11111111_11111110_00010011_01110110_11011010_11111111_11111111_00100000_01010101_10111100_10110110_11111111_11111111_11111111_10111011_11111111_11111111_11111111;
assign in[114] = 496'b11111111_11111111_11100010_01101001_01010010_11111111_11111111_11111111_11010101_01111101_00100010_11111111_11111111_11111111_11111110_00101101_01101010_11011010_11111111_11111111_11111110_00000010_01111101_10011000_11111111_11111111_11111111_10111111_01111101_01001101_11111101_11111111_11111111_11111101_00111101_01111101_10111110_11111111_11111111_11111111_11101011_01111101_01001110_11110111_11111111_11111111_11111111_10010110_01111101_10001100_11111111_11111111_11111111_11101100_01100001_01001110_11110011_11111111_11111111_11000000_11111111_11111111;
assign in[115] = 496'b00101010_00100001_10110011_11000001_00010001_00100101_10001111_11111111_11111111_11111111_11101011_11110100_01100100_11111010_11111111_11111111_11111111_11111111_11110001_01010110_11111111_11111111_11111111_11111111_11111111_11111110_01000100_11001101_11111111_11111111_11111111_11111111_11111111_11011000_01000100_00000111_00011110_10111011_11111111_11111111_11111111_11110101_00100011_01000001_11100011_11111101_11111111_11101111_00100011_01111100_01000011_00110101_00100011_11011100_01001101_10010110_11110010_11111111_11111111_11111111_11111111_11111111;
assign in[116] = 496'b11111111_11111100_00011110_01111101_01111101_11111111_11111011_00101000_01101110_10011010_00011110_11111111_11100101_01000001_01001111_11100011_11111111_10010100_11111011_01011001_00110001_11111000_11111111_11110101_01100010_10111101_01111101_11010011_11111111_11111111_10010011_01111010_00000001_01011001_11111111_11111111_10011101_01110101_00011101_01000001_00001110_11111111_10110110_01111010_01001011_11101110_01101110_10111001_11100101_01011100_01100010_11101110_11111111_01111000_00100010_01111001_01000100_11010110_11111111_11111111_11111111_11111111;
assign in[117] = 496'b10001000_11010101_11011110_11101100_11111111_01110101_01000100_01100110_01111100_01100110_11001111_01110011_11100011_11111111_11111000_11010101_10001010_01011010_01011101_11011000_11111111_11111111_11111111_11110101_01110110_10110100_01100010_10011001_00101010_11001011_00001111_01111110_11111111_10111111_00110110_00110001_11001101_01101100_00110101_11111111_11111111_11111111_11001111_01100111_01010011_11101111_11111111_11111111_11110000_01001000_01101100_11100010_11111111_11111111_11111011_01001001_01110110_11000111_11111111_01111110_10101001_11111111;
assign in[118] = 496'b11100111_01000000_01110101_01101000_01101100_11000111_01011110_01000101_11011100_11111001_10111001_11100111_01100001_01000100_11110001_11111111_11111111_11111111_10111010_01111101_11000110_11110111_11111111_11110011_11111110_10101110_01111101_00101000_01101111_01010010_01111011_00010100_10101010_01111101_01111101_01111101_01110101_01000111_11000010_11010110_01111101_00110111_11000111_10010111_11101000_11111111_00111010_01110111_10100010_01010100_01111101_10010001_11111111_00110011_01111101_01111100_01111101_00101000_11100101_10010100_11010110_11100001;
assign in[119] = 496'b11111111_10100011_01110010_01110111_01101010_11111111_11011101_01110001_00010100_00110011_00111001_11111111_11111111_00100111_01001011_00010101_01100000_11101010_11111111_11111111_10010001_01111010_01111010_11001111_11111111_11111111_11111111_10111110_01110011_01111101_01001011_11110001_11111111_10000110_01111000_10101110_10101100_01111101_10101010_00001101_01101011_10111110_11111111_10101001_01111101_11100001_01111101_00000110_11011000_00010011_01101011_01001011_11111111_01111101_01110010_01110101_01011110_10001010_11111010_11001000_11110110_11111111;
assign in[120] = 496'b11111111_11101001_01111001_11100010_11111111_11111111_11111111_10111001_01000010_11111111_11111111_11111111_11111111_11111111_00110100_11000100_11111111_11111111_11111111_11111111_11001001_01000000_11111111_11111111_11111111_11111111_11111100_01000111_11010001_11110101_00000101_11111101_11111111_10101100_01011001_11111111_10011000_01110001_11111010_11111111_00111001_00110100_11101010_01100000_10101101_11111111_11110110_01111110_01111110_01111011_00111100_11111111_11111111_11111101_10100001_11101010_10010011_11101111_11111111_11111111_11111111_11111111;
assign in[121] = 496'b11111111_11110111_00001100_01111100_01001011_11111111_11111111_01010001_01111101_00000111_01010010_11111111_11111101_00100101_01010101_11111010_11111111_00010000_11111111_10111111_01111101_11001000_11111111_11110100_01001111_11111111_10111001_01111101_11110100_11111111_10000001_01110001_11111111_00011111_01111101_11100001_10010101_01101010_10101011_11000010_01111100_00111000_00010010_01111101_10001001_11111111_00001010_01111101_01101011_01110001_10010010_11111010_11111111_11110100_01110000_01111101_10100010_11111111_11111111_01011000_11111010_11111111;
assign in[122] = 496'b11111111_11100101_01101110_10010000_11111111_11111111_11111111_10001110_01111111_00011101_11111111_11111111_11111111_11111111_00100011_01111100_11000001_11111111_11111111_11111111_11111110_01100000_00110010_11111111_11111111_11111111_11111111_10101000_01111110_00010001_11111111_11111111_11111111_11111111_00100001_01110001_11100111_11111111_11111111_11111111_11110010_01110001_10000100_11111111_11111111_11111111_11111111_11110101_01101011_10111011_11111111_11111111_11111111_11111111_10010011_01111110_11011110_11111111_11111111_00111101_11110111_11111111;
assign in[123] = 496'b11111111_11111101_10010111_01011010_01110000_11111111_11111100_00111001_00111100_10111100_01110101_11111111_11111111_10100011_01011100_11110110_10011011_01011101_11111111_11110000_01100000_11000000_11111011_01010100_10100010_11111111_11100100_01011111_10110010_10011001_01000000_11111101_11111111_11111111_11010011_00100100_01111101_00100001_11111111_11111111_11111111_11111100_01000011_00100111_11101111_11111111_11111111_11111111_00011110_01001001_11110100_11111111_11111111_11100011_00110011_01011011_11010110_11111111_11111111_11110011_11111111_11111111;
assign in[124] = 496'b11111111_11111111_11111111_00000100_01111101_11111111_11111111_11111111_11111111_00110100_01010001_11111111_11111111_11111111_11111111_10010010_01111010_10101110_11111111_11111111_11111111_10010101_01111101_00001110_11111111_11111111_11111111_11011101_01101111_00011000_11110110_11111111_11111111_11111111_00101100_01100011_11111010_11111111_11111111_11111111_11011111_01111101_00101000_11111111_11111111_11111111_10011111_10111011_01101111_11011101_11111111_11111111_11111111_11001000_01011011_00100011_11111111_11111111_11111111_11000110_11111111_11111111;
assign in[125] = 496'b11111111_11111111_11111111_11111111_11111111_11110000_11111111_11111100_00110010_01111100_11100100_01111100_01101011_00101010_00111000_01111101_01111100_11100100_00011110_01110111_01111110_01111101_01111110_00000010_11111010_11111111_11110100_11100010_00010101_01111101_10111010_11111111_11111111_11111111_11111111_10011110_01111110_10111010_11111111_11111111_11111111_11111111_10111110_01111101_00001101_11111111_11111111_11111111_11111111_11101110_01101111_01011001_11110111_11111111_11111111_11111111_11111111_00110000_01111101_11111111_11111111_00001100;
assign in[126] = 496'b01000110_00000100_11100111_11111111_11111111_10111111_01101010_11111011_11111111_11111111_11111111_11111111_11110110_01101001_11011000_11111111_11111111_11111111_11111111_11111111_10100000_01011010_11100010_11111111_11111111_11111111_11111111_11111111_10010110_01101001_11010011_11111111_11111111_11111111_11111111_11111011_00101100_00010100_10101010_11111111_11111111_11010011_00110110_10101111_11111011_00001001_11111111_11111111_01011010_11100111_11111011_10010110_01001011_11111111_11111111_00000100_01100100_01001011_00000100_11111111_11111111_11111111;
assign in[127] = 496'b11111111_11111111_11111111_11111111_11111111_11011111_10111110_00001111_10100010_11010110_11111111_01000101_00011110_00011110_01100111_00010000_01011010_00110100_11111101_11111111_11111100_00111011_11100011_11111100_00000101_11111111_11111111_11101001_01011111_11111111_11111111_11111111_11110111_11111111_10100001_00001000_11111111_11111111_11111111_00100101_11001110_01001100_11011101_11111111_11111111_11111111_10110011_10000011_11000110_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111;
assign in[128] = 496'b11111111_11111111_11111111_11111111_11111111_10000010_01001100_01111110_00110110_11000100_11111111_00001100_01001001_11001111_10111111_00111111_01111100_11000000_01001100_11110001_11111111_11111111_00110111_01111110_01000000_00110000_11111111_11111101_10001000_01111001_10100100_01011001_01011100_00101000_01010001_01100101_11000011_11111111_01001111_11000111_00101101_10000001_11110110_11111111_11111111_01011001_11111111_11111111_11111111_11111111_11111111_11011101_01011110_11111111_11111111_11111111_11111111_11111111_00001110_11111111_11111111_00000111;
assign in[129] = 496'b11111111_10101010_01111001_11010000_11111111_11111111_11111100_01100001_00100011_11111111_11111111_11111111_11111111_10010010_01111101_11011010_11111111_11111111_11111111_11111011_01011000_00011000_11111111_10011101_11001000_11111111_10010010_01111011_11110010_10110001_01111110_00000110_11111010_01011111_00010010_11111111_00111011_01111001_11010001_10011001_01111110_01000100_01001100_01111110_01001000_11111111_00000011_01111110_01111110_01101110_01010000_11001010_11111111_11101011_10000110_11001011_11111111_11111111_11111111_11111111_11111111_11111111;
assign in[130] = 496'b10000011_00111101_11111111_11111111_11111111_11111111_10111101_01111000_11100110_11111111_11111111_11111111_11111111_11101100_01111111_10110000_11111111_11111111_11111111_11111111_11101100_01111110_10110000_11111111_11111111_11111111_11111111_11101100_01111111_10110000_11111111_11111111_11111111_11111111_11110000_01111000_10110000_11111111_11111111_11111111_11111111_11111111_00111011_10000101_11111111_11111111_11111111_11111111_11111111_10000100_00001011_11111111_11111111_11111111_11111111_11111111_10011111_00001011_11111111_11111111_10101100_10011110;
assign in[131] = 496'b11110010_01100110_11001100_11111111_11111111_11111111_10100010_01001011_11111111_11111111_11111111_11111111_11111110_01100000_10011100_11010001_11111101_11111111_11111111_10101000_01111110_01111110_01111110_01010110_10110100_10111100_01111101_01100000_11000110_11101110_01011110_00111101_00110001_01111101_10000010_11111111_11111111_01010101_01011011_00001110_01011101_11111001_11111111_11110110_01011010_10001000_11011111_01101110_10001001_10101111_01001010_01010110_11110010_11111111_10111010_01000101_01110111_01000001_11100110_11111111_11111111_11111111;
assign in[132] = 496'b10000011_00010100_11010000_10110101_00011011_10100111_10001000_11111111_11111111_11111111_10011011_11111011_00110000_11111100_11111111_11111111_11111111_11010011_11000111_10010011_11111111_11111111_11111111_11111111_11010111_10101100_10110010_11111111_11111111_11111111_11111111_11001011_10101100_10110010_11111111_11111111_11111111_11111111_10010000_11000000_10101000_11111111_11111111_11111111_11111010_00101100_11110000_00001101_11111111_11111111_11111101_00000000_10111110_11111111_00011100_11110110_00010101_01011110_10000100_10000001_10001001_11110001;
assign in[133] = 496'b11111111_00011110_10001010_11111111_11111111_11111111_11111111_01100101_11100100_11111111_11111111_11111111_11111111_10101001_00001010_11111111_11111111_10110110_11111111_11000011_01011010_11100001_11111111_11011100_01100010_11101000_01100000_01111110_01101101_01011101_01101011_00010101_11111111_00001110_10110011_10101001_01111000_00000111_11111111_11110111_00110011_11111111_11111111_01001010_11100011_11111111_10000001_10100011_11111111_11111111_00001110_11110101_11111111_01101101_11011100_11111111_11111111_11111111_11111111_11111111_11111111_11111111;
assign in[134] = 496'b11111111_11111111_11111111_11111111_11111111_11111111_10110101_01010100_01101001_00011111_11101111_11111111_11100010_01100110_01010100_01110000_01011111_01000111_11111111_00111110_10101010_01001110_10100101_11101000_01010101_11001000_01011111_00011111_01001101_11111100_11111111_00100111_10110100_01111110_01010011_11100010_11111111_10110001_00100010_11101110_00001110_11010100_11111111_11100010_00110000_11010001_11111111_11111111_11111111_11111100_00111101_10101000_11111111_11111111_11111111_11111111_00100100_00011011_11111011_11100001_01001100_11110100;
assign in[135] = 496'b01111010_11000001_11111111_11110110_10000100_11101111_01011010_00011101_11100100_01010011_01001111_11111111_11111111_10001011_01111110_01101101_01101101_00011110_11111111_11111111_11011101_01110011_00110101_10000111_10001011_11111111_11110111_01010011_10000110_11111111_11111111_11111111_11110100_00111101_01001001_11111001_11111000_11111100_11111111_00010001_01111110_00001101_10100010_01110100_00100000_11111111_01001110_00110001_11101011_01100101_01100110_11100011_11111111_01110011_01110110_01101110_01101100_11001011_11111111_01000101_00000001_11111111;
assign in[136] = 496'b10100000_11111111_11111111_11111111_10110100_01101001_01011010_11111111_11101100_00111100_01111101_11111111_10010110_01111000_10010000_01010000_01111001_01101110_11111111_11101100_01011010_01111101_01111101_01111101_01010101_11111111_10110100_01101001_01011111_00001001_11000011_11111111_10111001_01111000_00101101_11010011_00110110_10111001_11111111_01000110_01010110_11001110_01011111_01111101_10100000_11111111_01111110_00001110_01010101_01111101_01000110_11110110_11111111_01111110_01110100_01111101_01000001_11111011_11111111_10100000_11111011_11111111;
assign in[137] = 496'b11111111_11101110_01010111_10000101_11111111_11111111_11111111_10000010_01010100_11111110_11111111_11111111_11111111_11110100_01101111_10110110_11111111_11110011_11111111_11111111_00011000_01000011_11111111_11011001_01110010_11111111_11101011_01110010_10110000_11111101_01010011_01101101_11111111_10000011_01111110_11011001_10101000_01111110_10010100_11011101_01110010_01010011_10011000_01101100_00101001_11111111_10101001_01111110_01111110_01111110_01100000_11110110_11111111_11111011_10011011_11010111_11001011_11111010_11111111_11111111_11111111_11111111;
assign in[138] = 496'b11111111_11111111_11111111_11111111_11000000_00010100_11010110_11111100_10100100_01001010_01111101_11001000_01111010_01110111_01001011_01111101_01011000_01111101_11111111_11011111_01000001_01111100_01111101_01111100_01001011_11111111_10010010_01111001_01000100_00101011_11000000_11111111_11010101_01101110_10001110_11111111_10011001_10100110_11111111_00011100_00100000_11111111_11011111_01110010_10011100_11111111_01111000_10011100_11100001_01001010_01011110_11101010_11111111_01111110_10011000_01011101_01110010_11000000_11111111_00111010_11011000_11111111;
assign in[139] = 496'b11111111_10000100_01101101_11100001_11111111_11111111_11011110_01101001_00110101_11111111_11111111_11111111_11111111_00100001_01111101_11000101_11111111_11111111_11111111_11011011_01111100_00101110_11001010_00101110_01001001_11111111_00110000_01111110_01110001_01111111_01111110_01111010_11000011_01111101_01111110_01000011_00010011_01111100_00010010_10111100_01111110_01010011_00111010_01111000_01001111_11101000_10111001_01111110_01111110_01101001_10010111_11110110_11111111_11101101_01001100_00010101_11011100_11111111_11111111_11111111_11111111_11111111;
assign in[140] = 496'b11111000_10001111_01011000_01111101_01110001_11111111_00001011_01111100_01001011_00110100_01000011_11111111_10100100_01111100_10011011_11111111_11111111_11101100_10110111_01110011_10001011_11111111_11111111_11111111_00101000_01110101_00001010_11111111_11111111_11111111_10110110_01111011_01111101_11001110_11111111_11111111_11110010_01010000_01100001_01111101_11000100_11111111_11110001_00100100_01110110_10110111_01111101_00110101_11101010_00110010_01111101_10001110_11111111_01111101_01111101_01001000_01101111_10101000_11111111_01111000_10100011_11111111;
assign in[141] = 496'b10110110_00110110_01011010_01001010_11001000_10011000_01010000_10111110_11111001_10011100_01100000_11000001_01000110_11111010_11111111_11111111_11110110_01111101_00011000_10110111_11111111_11111111_11111111_11111001_01110011_00010111_11110111_11111111_11111111_11111111_10110111_01100010_01000101_11111111_11111111_11111111_11111101_01000100_10011010_01010111_11111111_11111111_11111111_10010001_01001010_11111101_00000100_00011101_00101010_11010101_01101011_11001110_11111111_11111111_01011000_11000100_01001111_10101001_11111111_01101101_10110100_11111111;
assign in[142] = 496'b11111111_11111111_00111000_10000101_11111111_11111111_11111111_10111011_01011110_11110011_11111111_11111111_11111111_11111111_00111110_10010110_11111111_11111111_11111111_11111111_10011100_01111101_10010100_11111110_11111111_11111111_11101000_01110000_01000011_01100000_01100000_11011000_11111111_00101011_01000011_11111011_11111111_01011011_10011100_11100110_01111110_11001000_11111111_11001110_01101101_11001010_11111001_01101000_00111001_00111001_01111001_00011100_11111111_11111111_11100101_10010001_10000001_11001110_11111111_11111111_11111111_11111111;
assign in[143] = 496'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11110101_10110011_10001100_10100001_10100001_00100000_00111010_01101110_01111101_01111101_00110011_00110011_00010111_10010010_10001111_01111100_01001010_11111111_11111111_11111111_10100101_01110000_10000101_11101001_11111111_11111111_10010110_01101101_10101111_11111111_11111111_11111111_11101111_01101011_10111000_11111111_11111111_11111111_11111111_11001010_01111101_11011110_11111111_11111111_11111111_11111111_11001010_01110100_11100111_11111111_11111111_01000010_00010100_00110001;
assign in[144] = 496'b11111111_11111111_11111111_11111111_11110000_01111101_10101100_11111111_11111111_10101011_01110011_11111111_00101010_01001000_11010110_00010100_01111100_01010010_11111111_00001010_01111101_01111101_01111101_01100101_01011001_11111111_11111100_00111000_01101110_01000000_01000000_00111010_11111111_10010100_01111011_00010111_11111111_11111111_11111111_10001001_01110111_00001100_11111001_11111111_11111111_11111111_01110011_00010100_11111111_11111111_10100110_11101011_11111111_01111101_11001100_11111111_00001111_01111101_10101101_01001010_01100100_10101000;
assign in[145] = 496'b11110100_01111010_00011011_11111111_11111111_11111111_11110011_01111110_00011011_11111111_11111111_11111111_11111111_11110011_01111101_00011011_11111111_11111111_11111111_11111111_11110011_01111101_00011011_11111111_11111111_11111111_11111111_11110011_01111110_10011100_11111111_11111111_11111111_11111111_11011000_01111101_11001011_11111111_11111111_11111111_11111111_10101100_01111110_00011011_11111111_11111111_11111111_11111111_10111000_01111101_00011011_11111111_11111111_11111111_11111111_11110011_01111101_10000001_11111111_11111101_10010001_11111001;
assign in[146] = 496'b10000011_10000001_00001111_01000111_10111010_01011001_01100001_00010110_00010000_01110100_10001110_11000111_01111100_11100101_11111111_11111111_11111111_11111111_10111010_01111101_11100101_11111111_11111111_11111111_11111111_11111010_01011111_01010001_00000011_10000011_10110000_11111111_11111111_11100110_00101001_01111101_01111101_01010011_11111111_11111111_11111111_11111111_11111111_10001111_01010011_11111111_11111111_11111111_11111111_11111111_00011000_01010011_11111111_11111111_11101111_11100001_00010101_01111101_00101101_01111110_00111000_10101011;
assign in[147] = 496'b11111111_11111111_11111111_11111111_11111111_11111111_11010111_10010011_00011010_00111011_01111110_11111111_10011110_01111000_01111010_01101000_01111110_01111110_11100001_01101001_10011100_11010001_01101000_00001001_01011111_10001111_00111010_11111011_01010001_00111011_10010000_01011010_00011111_00010000_10010101_01011111_01000000_01101011_11100011_10011010_01110111_00101010_10100100_01111100_00011001_11111111_11111111_11000101_11111010_00010100_01111010_11001110_11111111_11111111_11111111_11101110_01111100_00000101_11111111_00111001_01011110_11101010;
assign in[148] = 496'b01101111_10001111_11111111_11111111_11111111_11111111_00101000_10010000_11111111_11111111_11111111_11111111_11111111_00111111_10010000_11111111_11111111_11111111_11111111_11100100_01110110_10011111_11111111_11100001_11111111_11111111_11000001_01101010_11001000_00110011_01110110_01011111_11111111_10000010_01111000_01110110_00101011_11000011_01111110_11111110_01001110_01111100_10011011_11111001_10010001_01011001_11110111_01100000_00110100_00111100_01010001_01101101_11010011_11111111_11111111_11111111_10101010_10100001_11111010_11111111_11111111_11111111;
assign in[149] = 496'b11111111_11011101_10000010_10101010_11111111_11111111_10111110_01100000_00001001_01111110_11100111_11111111_11110001_01100100_11011101_11111111_01010000_11001101_11111111_11010010_01011010_11111111_11100111_01111000_11011101_11111111_11111111_00100111_00010011_01010000_01000110_11111111_11111111_11111111_11111111_11101100_01011010_11000011_11111111_11111111_11111111_11111111_10011011_00111100_11111111_11111111_11111111_11111111_11111011_01011111_11000011_11111111_11111111_11111111_11111111_10010001_00110010_11111111_11111111_01100100_11101100_11111111;
assign in[150] = 496'b11111111_11111111_11000101_01011001_01111100_10011001_10001000_10011001_01101111_01111100_01111100_11111111_01001111_01111100_01111101_01111100_01111100_01111100_11111111_10011011_01111100_01111101_01111100_01111100_01111100_11111111_01001111_01111101_01111110_01111101_01111101_01111001_10111101_01111100_01101010_10010111_00010101_00000011_11100110_00101100_01111100_00111111_11111111_11111111_11111111_11111111_00110101_01111100_00101111_10100111_10110000_11111110_11111111_10001000_01111100_01111100_01111101_01110111_11011011_01111101_01100111_10100100;
assign in[151] = 496'b11111111_11110000_00100100_01111100_01111101_11111111_11100011_01010101_01110110_10001110_11011000_11111111_11101011_01010111_01110101_10111111_11111111_11111111_11111111_10110100_01111101_00111010_10100010_11111110_11111111_11111111_11011110_01011001_01111101_01111101_11111000_11111111_11111111_11111111_00010110_01111101_00001010_11111110_11111111_11111111_11101101_01110001_00101001_11111111_11111101_11111111_11111111_11011000_01111101_10110101_00011111_01010111_11110001_11111111_11011000_01111101_01111100_01110000_00010101_10010010_10001110_11011111;
assign in[152] = 496'b11111111_11010110_01011100_01101010_01001110_11111111_11011101_01101010_00101010_11111001_11001111_11111111_11111111_10001111_01000000_11111001_11111111_11111111_11111111_11111111_11101011_01010100_11010110_11111111_11111111_11111111_11111111_11111111_00000111_10010110_11111111_11111111_11111111_11111111_11111001_01011100_11000000_11111111_11111111_11111111_11111111_00010101_01001110_11111111_11111111_11111111_11111111_10011101_01101010_11001111_11000111_11111001_11111111_11100100_01111000_00010100_11000000_01101010_10111010_00000000_00000000_11000000;
assign in[153] = 496'b11010111_01111101_01111101_00110111_11111111_11111111_00110110_01111101_01111101_10111010_11111111_11111111_11010111_01111101_01111101_01010011_11111111_11111111_11110010_01100001_01111101_01111101_10111010_11111111_11111111_10111010_01111101_01111101_01010011_11111111_11111111_11111111_00110110_01111101_01111101_10111010_10101100_10000010_10000010_01010011_01111101_01101111_01010011_01111101_01111101_01111101_01010011_01111101_01111101_01111101_01111101_01111101_01010011_10000010_01111101_01010011_00011011_10101100_11110010_11111111_11111111_11111111;
assign in[154] = 496'b01011111_01111100_01111101_01111011_10011111_00100010_01111110_00100111_01010011_01111101_10000001_11111111_00001000_01111101_01000111_01111001_01110110_11000011_11111111_11101000_01100010_01111101_01111110_00110010_11111111_11111111_11111111_00011101_01111100_01111101_00101000_11111111_11111111_10111111_01110010_01111101_01111110_01111001_10110001_00100011_01110110_01111101_00001111_00010111_01111100_01000010_00100010_01111100_01111101_00100001_01100010_01111100_00100010_11000100_01011100_01111101_01111100_01111101_00100100_10000001_10000010_10111010;
assign in[155] = 496'b11111111_11111111_11111111_11111111_11111111_01001100_11111110_11111111_11111111_11111111_11100001_01011100_01111101_10011100_10100001_10100001_10000111_01100110_01111101_01111101_01111101_01111101_01111101_01111101_01111101_01111101_01111101_01111101_01111101_01111101_01111101_01111101_00101000_01111101_01011110_10100000_11110100_11110100_11000000_10000110_01111101_10010111_11111111_11111111_11111111_11100010_10011101_01111101_10111101_11111111_11111111_11111111_11100010_00010011_00100101_11111111_11111111_11111111_11111111_11111111_11111111_11111111;
assign in[156] = 496'b11111111_10111011_01011010_01100100_11010000_11111111_11001100_01111101_01111101_01111101_10111011_11111111_11111111_11010101_01101101_01111101_01111011_11001110_11111111_11111111_11010110_01111011_01111101_01000011_11111111_11111111_11111111_10100101_01111101_01111101_10010001_11111111_11111111_11111111_00000110_01111101_01111101_10100100_11111111_11111111_11010101_01110110_01111101_01100111_11011010_11111111_11111111_11000100_01111100_01111101_10001101_11111111_11111111_11111111_11001000_01111100_01110101_10111100_11111111_01100000_00101001_11111111;
assign in[157] = 496'b11111111_11110010_10001101_01010110_01111100_11111111_11010001_01100101_01111100_01101100_01101110_00011100_00011111_01100110_01111101_00100011_11011000_01010011_00100001_01111100_01111100_01111101_10100011_01100010_01111100_11011001_01111101_01111101_01111110_01111101_01111101_00111011_11011001_01111100_00111111_11001100_10111110_11011010_11111111_11011111_01111000_01100000_11101010_11111000_11011111_11111111_11111111_00011111_01111100_01101000_01100111_01101110_11101111_11111111_10001111_01111100_01111101_01100101_00000111_01000010_10111100_11110010;
assign in[158] = 496'b11111111_11111101_11010011_10010100_11010001_11111101_10001011_01011011_01111100_01110000_01100001_11011001_00110100_01100101_10111001_10100011_01111110_01001100_00001011_01110010_11000010_10010001_01101111_01100100_00101101_01000100_01111100_01110100_00110000_11001011_00011000_00111001_11100001_10111011_11100010_11111111_11010000_01100010_10000010_11111111_11111111_11111111_11110010_01010010_00111111_11111111_11111111_11111111_11101001_00100011_01100000_11100001_11111111_11111111_10011110_01100111_00100001_11011110_11111111_10000101_11111111_11111111;
assign in[159] = 496'b11111111_11111111_11111111_11111111_11111111_10011110_01111110_01111101_00001111_11111111_11111111_00100011_00010111_11110011_11100101_01001100_00111111_11101111_00000101_11000110_11100110_10110101_01000100_01111101_11011000_10100110_01110011_01010001_00101110_10100001_01101111_11011000_11111011_10100111_11110101_11111111_11000111_01110000_11101101_11111111_11111111_11111111_11111111_10010110_01000100_11111111_11111111_11111111_11111111_11111111_00000111_10001101_11111111_11111111_11111111_11111111_11101101_01011100_10111011_11111111_11000100_01100011;
assign in[160] = 496'b11111111_11110011_00100010_01111101_01001110_11111111_11111111_11010101_01111101_01111101_01101100_11111111_11111111_11111111_10001101_01111101_01111101_10011000_11111111_11111111_10111111_01111010_01111101_01100110_11111010_11111111_11111111_00111000_01111101_01111101_00001001_11111111_11111111_11001110_01111001_01111101_01101101_11100101_11111111_11111111_10011100_01111101_01111101_10010001_11111111_11111111_11111111_01010110_01111101_01011101_11110110_11111111_11111111_11111111_01101100_01111101_00010001_11111111_11111111_01011010_11110101_11111111;
assign in[161] = 496'b11111111_11111111_11111111_11101010_11010000_11111111_11111100_10100001_00110111_01110011_01111101_11110110_10110101_01000111_01111101_01111011_00100101_01001111_01110110_01111101_01111101_01111101_01011001_00101110_01111001_01011110_01111101_01110100_01111101_01111101_01111101_01100111_01011110_01111101_10101100_11011110_11011110_11011110_11110101_01110111_01011010_11111111_11111111_11111111_10110101_10000111_01011101_01111101_00010101_00101100_01101011_01111101_01111101_10111101_01110100_01111101_01111101_01111000_01001001_11010000_11010000_11011110;
assign in[162] = 496'b11101110_01111110_11101101_11111111_11111111_11111111_11011000_01110000_11111111_11111111_11111111_11111111_11111111_10101110_01001101_11111111_11111111_11111111_11111111_11111111_10010100_00100011_11011000_11111111_11111111_11111111_11111111_00011111_01111110_01111101_00000110_11111111_11111111_11111111_01101001_00101101_11001101_01110011_11110111_11111111_10111110_01110101_11110010_11111000_01101001_10011110_11111111_11110000_01011010_10101111_10010011_01110010_11101010_11111111_11111111_10111110_01101100_01000100_10111000_11111111_11111111_11111111;
assign in[163] = 496'b11111111_11100011_01100101_01111101_01011001_11111111_11111000_01000010_01111110_01110111_10110101_11111111_11100010_01011000_01111101_01110101_10110100_11111111_11111111_00110010_01111110_01111110_10100011_11111111_11111111_11000101_01111101_01111101_00010100_11111111_11111111_11111111_01011000_01111101_01111101_10110001_10011111_10010011_10101111_01111101_01111101_01111101_01111101_01111110_01111101_01111101_01101100_01111101_01111101_01111101_01011011_00111001_10110000_11101110_10101011_10011000_11001010_11111010_11111111_11111111_11111111_11111111;
assign in[164] = 496'b01111100_01111101_01111100_01111100_01011100_01111100_01111100_00111010_01011101_01111100_01011111_11011011_01111100_01111100_00110011_01111001_01111100_10101111_11011011_01111100_01111100_01111101_01111100_00000101_11111111_11011011_01111101_01111101_01111110_01001010_11111111_11111111_01010101_01111100_01111100_01111101_01111100_10010010_11111111_01111100_01011111_00000111_10001001_01101110_01111100_10101111_01111100_01110010_00001111_10001001_01010001_01111100_01110010_10000001_01111001_01111100_01111101_01111100_01111100_10000010_10000001_10000010;
assign in[165] = 496'b10010001_00100001_11011110_11101001_11111111_11000101_01101011_11100110_11111111_11111111_11111111_11111111_00110010_10010100_11111111_11111111_11111111_11111111_10110101_01011100_11111011_11111111_11111111_11111111_11111111_10111011_01011110_01011110_00101001_10001111_11101011_11111111_11111111_11111011_10111001_10110010_00010111_01100100_10100001_11111111_11111111_11111111_11111111_11111111_10100011_00010100_11111111_11111111_11111111_11111111_11100000_01010000_10111110_11111111_11110101_10110011_00011001_01010110_10110001_10000011_11000001_11110101;
assign in[166] = 496'b11010111_10001011_10111010_11111111_11111111_00010000_01110010_01011000_01111000_11000010_11111111_10100010_00011101_11101101_11111100_01100011_01110000_11011110_01000001_11111001_11111111_10010010_00100011_00101110_10111100_10000001_11111010_10001111_00111111_11101011_10000010_10100000_01100001_01100110_00010110_11110101_11111111_00001110_10010001_11110010_11101111_11111111_11111111_11111111_01001010_10101111_11111111_11111111_11111111_11111111_11101100_01101100_11100101_11111111_11111111_11110011_11111111_00001100_00001110_10111110_00010110_01001101;
assign in[167] = 496'b11111111_11100001_01000010_01111001_11001100_11111111_11111111_01000011_01111100_01111100_10011001_11111111_11111111_11111111_01010011_01111101_01100111_11100100_11111111_11111111_11000011_01111010_01111100_00001101_11111111_11111111_11111111_00101000_01111110_01110001_11001100_11111111_11111111_11111111_01101110_01111101_00100000_11111111_11111111_11111111_11111111_01101110_01111101_10001011_11111111_11111111_11111111_11111111_01101111_01111110_11110001_11111111_11111111_11111111_11001100_01111100_01001110_11111111_11111111_01110001_00100100_11111111;
assign in[168] = 496'b10000010_00101011_00101011_00101011_10011111_01101010_01111101_01111101_01111101_01111101_01111101_01111101_01111101_01101011_00111110_00010100_00010100_01101011_01111101_00100001_11110011_11111111_11111111_11111111_00010011_01111101_10111111_11111111_11111111_11111111_11111111_01010100_01111101_00110101_11100101_11111111_11111111_10100110_01111001_01111101_01111101_01100100_10111000_11011010_01011001_01111101_01111101_01111101_01111101_01111101_01110101_01111101_01111101_10010110_01101010_01111101_01111101_01111101_01101101_10110000_10001110_00101100;
assign in[169] = 496'b11111010_00100010_01010011_00110111_10110100_11111111_00000110_10010011_11111111_11111111_00010100_11111111_11111111_01000101_11110110_11111111_11111111_11110100_11111111_11111111_00111000_11111111_11111111_11111111_11111111_11111111_11111111_00101101_11001111_10010100_10001111_11111111_11111111_11111111_11100000_01101110_01100101_10000100_11111111_11111111_11111111_10101010_00001111_11111111_11111111_11111111_11111111_11111111_01001001_11100111_11111111_11111111_11111111_11111111_11111111_01011001_11110000_10101110_11111111_10100100_01010111_01100000;
assign in[170] = 496'b11111111_11110000_00001011_01011001_11000101_11110100_10001111_01101000_01110100_10000011_11111110_10110100_01010000_01111010_00111000_11001111_11111111_11111111_01111110_01010001_11010011_11111111_11111111_11111111_11111111_01111111_00000011_11111111_11111111_11111111_11111111_11111111_00110010_01101001_00001101_11011111_11111111_11111111_11111111_11111010_00101000_01101001_01111010_00111001_10001000_10010100_11111111_11111111_11110100_10000010_01010001_01111110_01111110_11111111_11111111_11111111_11111111_11111101_11101001_11111111_11111111_11111111;
assign in[171] = 496'b11111111_00001100_01111100_01001011_11111111_11111111_11100011_01111001_01111010_10100000_11111111_11111111_11111111_01000010_01111101_00000001_11111111_11111111_11111111_10101101_01111100_01011101_11110001_11111111_11111111_11110001_01011111_01111100_01111101_01011011_00111001_10111101_11011101_01101110_01111100_00111001_00101001_01101110_01100111_11100101_01010010_10100100_11111111_10111111_01101100_00111100_00100001_00100101_10010100_00110111_01110111_01100100_11010101_00010010_01011001_01111101_01101110_00001101_11101110_11111111_11111111_11111111;
assign in[172] = 496'b11111111_10111001_01010110_11100001_11111111_11111111_11111111_11000100_01111101_11011001_11111111_11111111_11111111_11111111_11000110_01111101_11011101_11111111_11111111_11111111_11111111_00000101_01100011_11111111_11111111_11111111_11111111_11111111_00010011_01000011_11111111_11111111_11111111_11111111_11111111_00111010_00010011_11111111_11111111_11111111_11111111_11111111_01101100_00001111_11111111_11111111_11111111_11111111_11011110_01111101_10101101_11111111_11111111_11111111_11111111_11011001_01111110_11100000_11111111_11101000_01011110_11110111;
assign in[173] = 496'b10010001_01000000_01111111_01101111_01000000_01100000_01111111_01111111_01111111_01111111_01111111_00110000_01111111_01010000_11000000_11111111_11111111_00100000_01111111_01111111_10110000_11111111_11111111_11111111_10100000_00010000_01111111_01010000_00000000_11000000_11000000_11110000_11111111_00000000_01111111_01111111_01111111_01111111_10010001_11111111_11111111_00101111_01111111_01101111_00100000_11110000_11111111_10010000_01111111_01000000_11110000_11100000_11000000_11111111_01000000_01111111_01010000_01101111_01111111_01000000_01111111_01111111;
assign in[174] = 496'b11111111_11111111_11101000_10111011_11001101_11111101_10100010_01011001_01111101_01101110_01011010_11111111_10110010_01111110_00111010_10111011_11111111_11101011_11111111_00011111_01111110_11001111_11111111_11111111_11111101_11111111_11110011_00100110_01100011_10000110_11111000_11111111_11111111_11111111_11110011_00100001_01111110_01110000_10011000_11010101_10100011_00000000_00101010_01111001_00101010_11110010_01111110_01111110_01111001_00110101_10100110_11111001_11111111_11000101_11010000_11100111_11111111_11111111_11111111_11111111_11111111_11111111;
assign in[175] = 496'b11111111_11111111_11111111_11111111_11111111_10000111_00100010_10111100_11111101_11111111_11111111_11111111_11111111_11110000_10001110_01010110_00111110_00011101_11111111_11111111_11111111_10010011_10100001_11100011_00010100_11111111_11111111_10110100_10001001_11111111_11111111_11111111_11111111_11111110_00100111_11111001_11111111_11111111_11111111_11111111_11010111_10100001_11111111_11111111_11111111_11111111_11111111_10101001_10111100_11111111_11111111_11111111_11111111_11111111_10101001_10111010_11111111_11111111_11111111_00011110_11010100_11111000;
assign in[176] = 496'b11111111_10001001_01111100_01101011_11100011_11111111_11001010_01110100_01111010_10110001_11111111_11111111_11111111_01100110_01111101_00101000_11111111_11111111_11111111_10001100_01111101_01101010_11100101_11111111_11111111_11001000_01110110_01111001_10110101_11111111_11111111_11111111_00110100_01111100_10001000_11111111_11111111_11111111_11001110_01111100_01110011_11001011_10011011_00011001_01011110_01111001_01111100_01111100_01111100_01111101_01111100_01110000_01011010_10100001_10111110_10000110_10111100_11000010_11111100_11111111_11111111_11111111;
assign in[177] = 496'b11111001_01000111_00111110_00001110_00110011_11111111_10110011_01010100_11111010_11111111_11111111_11111111_11111111_10101100_01110111_11100100_11111111_11111111_11111111_11111111_11110101_01010011_00010101_11111111_11111111_11111111_11111111_11111111_11001011_01101110_10101111_11111111_11111111_11111111_11111111_11111111_00101010_00010010_11111111_01101000_00110000_11001000_11000011_00110100_00000110_11111111_10101111_00100100_01111101_01111101_01001001_11110110_11111111_11001110_00100010_01111101_00111010_11110110_11111111_10101100_11111111_11111111;
assign in[178] = 496'b11110011_10101100_10100110_10100111_11011111_10000010_01110010_01111101_01111110_01111101_01111101_01100100_01111100_01111101_01110110_01010111_01010110_01111001_01111110_00011000_11001010_11011101_11111111_11111111_01000110_01111101_11101110_11111111_11111111_11111111_11110000_01101001_01111110_11011111_11111111_11111111_11111111_00010011_01111101_01111101_01110000_00110001_00001000_10000010_01110001_01111100_01110001_01111100_01111101_01111100_01111101_01111100_00101110_11110010_10101011_10100101_10100001_00100011_10010001_11111111_11111111_11111111;
assign in[179] = 496'b11111111_11111111_01000101_11000011_11111111_11111111_11111111_11011010_01011100_11111111_11111111_11111111_11111111_11111111_10001011_00100001_11111111_11111111_11111111_11111111_11111111_01010001_10111011_11111111_11111111_11111111_11111111_11111111_01111011_11011010_11111111_11111111_11111111_11111111_10110001_01011101_11111111_11111111_11111111_11111111_11111111_00011111_00010100_11111111_11111111_11111111_11111111_11111101_01100110_11010010_11111111_11111111_11111111_11111111_11010110_01111001_11111110_11111111_11111111_10101100_11111111_11111111;
assign in[180] = 496'b11111111_11111111_11101110_10100010_11111001_11111110_11111111_11011110_01010010_01111101_10010110_11000100_01001100_00111100_01011101_01011000_00010101_10010000_11100101_10111001_00100010_01111110_01011001_01010101_10100100_11111111_11111111_01001000_00111110_00000000_10100101_11111111_11111111_11111111_01110110_10111100_11111111_11111111_11111111_11111111_11111111_01110110_11001100_11111111_11111111_11111111_11111111_11111111_01110110_10101010_11111111_11111111_11111111_11111111_11111111_00100010_01001101_11111010_11111111_11110000_01100100_01011110;
assign in[181] = 496'b11111111_11111111_11111111_11111111_11111111_10010000_11111111_11111111_11111111_10110000_00110000_11111111_00101111_00110000_10110000_00101111_10010001_11111111_11111111_11111111_00100000_01111111_01100000_00000000_00010000_11111111_11010001_01100000_11010001_11111111_11010000_11111111_11111111_01000000_11010001_11111111_11111111_11111111_11111111_11100000_01101111_11111111_11111111_11111111_11111111_11000000_00000000_00000000_11111111_11111111_11010000_00010000_00000000_10010001_00101111_10110000_00100000_01000000_11010001_10110000_11010000_11111111;
assign in[182] = 496'b11111111_11100110_01110010_00011111_11111111_11111111_11111111_00011100_01111101_10000110_11111111_11111111_11111111_10110010_01111100_01000101_11111111_11111111_11111111_11001101_01110010_01111101_00011111_11001101_11110010_11111111_01000100_01111101_01011100_01101111_01111100_01111101_11010010_01111101_01001111_11111101_11010111_01111101_01111101_01010110_01110010_11011001_11111111_00010011_01111000_10011101_01111110_10001111_11111111_11111010_01000000_10011100_11111111_00100011_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111;
assign in[183] = 496'b00001001_00000101_00100111_00010001_11111111_11111111_11111010_11111111_10111010_01111011_11110011_11111111_11111111_11111111_11111111_10011000_01010000_11111110_11111111_11000111_10001110_10000010_01010111_00110011_10111010_11011001_01001101_00011011_01010110_01100010_00011011_01010010_11111111_11111011_11010111_01101100_11010000_11111111_11111111_11111111_11110000_01010010_10001000_11111111_11111111_11111111_11100111_00110010_01001000_11111110_11111111_11111111_11111111_01101100_01100011_01010011_00111100_11000010_11111111_11111100_11000111_10100100;
assign in[184] = 496'b11111111_11111111_11111111_11111111_11111111_00001001_00110001_01010101_01111100_00110110_10011000_01111101_01101100_01001111_01001010_01100100_01111101_01111100_01011100_11001001_11001110_10110111_01001111_01111110_01111101_01111101_01111100_01111101_01111100_01100111_01111011_01111100_11011001_10111010_11001010_11000010_10110001_01111010_00111111_11111111_11111111_11111111_11100010_01010011_01110111_10111100_11111111_11111111_11111111_00111110_01111100_10000001_11111111_11111111_11111111_10101010_01111101_00110000_11111101_01101001_01011010_11100111;
assign in[185] = 496'b11111111_11111111_01000000_10110100_11111111_11111111_11111111_11010111_01001100_11111101_11111111_11111111_11111111_11111111_00100000_10110010_11111111_11111111_11111111_11111111_11001001_00110010_11111111_11111111_11111111_11111111_11111111_00111000_10101000_11111111_11111111_11111111_11111111_10110111_01111110_11101110_11111111_11111111_11111111_11111111_00011101_01000011_11100110_11111011_11111110_11011101_11111111_00100010_01111000_01110110_01100000_00110110_01001000_11111111_11100011_10001110_11011010_11111111_11111111_11111111_11111111_11111111;
assign in[186] = 496'b11111111_01111001_00001110_00111101_01000110_11111111_11111111_01101001_11111000_00011111_00111111_11111111_11111111_11111111_01100110_11101000_01011111_10111100_11111111_11111111_11111111_01101011_01100001_01011101_11101101_11111111_11111111_11100100_01101011_01111100_10110100_11111111_11110010_10001100_01101000_01000000_00111111_00011001_11111010_01011101_01011001_10100110_11111001_11101011_01100101_11011000_01111011_00011000_10110001_11100101_10100110_01011110_11100101_10111000_00110000_01110000_01011110_00111011_10001101_11111111_11111111_11111111;
assign in[187] = 496'b11111111_11111111_11111111_11111111_11111111_10101100_01000101_01111110_01111110_01111110_01001001_01100000_01111110_01111110_01111110_01110000_01111000_01111110_01111110_01111110_01001110_00110100_10100001_01100010_01111110_01111110_01111110_01111110_01111110_01111110_01111110_01111110_01010100_01011101_01011101_01000100_01010000_01111110_01111110_11111111_11111111_11111111_11111111_01001011_01111110_01001011_11111111_11111111_11111111_10001111_01111110_01100100_11101001_11111111_11111111_10111000_01110101_01111110_10110010_01110101_01111110_00110100;
assign in[188] = 496'b11111111_11111111_11110110_10011011_11111111_00000100_11101100_11111111_00011000_01111101_11101100_00001110_01010101_01110011_10100101_01110011_00011000_11111111_11111111_11110110_01001011_01111101_01011111_11111111_11111111_11111111_11111111_11000011_01111101_00101100_11111111_11111111_11111111_11111111_11100010_01111101_11000011_11111111_11111111_11111111_11111111_10011011_01111101_11111111_11111111_10111001_11111111_11111111_10101111_01111101_11011000_10101111_01110011_11111111_11111111_11110110_01011111_01101001_01110011_11111111_11101100_10111001;
assign in[189] = 496'b00010110_01111011_01111110_01000110_01011011_10100010_01111000_00000110_11100000_11111111_11111111_11111111_01001010_00000100_11111111_11111111_11111111_11111111_11111111_00110000_10000101_11111111_11111111_11111111_11111111_11111111_11110000_01001010_00110010_11000100_11111111_11111111_11111111_11111111_10110110_01100010_01111000_11100110_11111111_11111111_10000110_01111101_00101101_10011011_11111101_11111111_11111000_01111000_00000101_11111111_11111111_11111111_11111111_11111111_00001111_01110101_01000101_00101011_00110010_11001101_10101110_10000001;
assign in[190] = 496'b11101111_01011100_01111010_11100010_11111111_11111111_10011110_01111101_00110111_11111111_11111111_11111111_11111110_01010101_01111101_10101110_11111111_11111111_11111111_11000010_01111101_01100001_10111100_11110110_11111111_11111001_00110111_01111101_01111101_01111101_01101101_01000101_00000010_01111101_01110101_00110000_00000000_00010111_01011011_10111100_01111001_01100001_10111110_11111111_11001101_01100010_11111111_11100000_01011110_01111011_00111000_01101100_00111110_11111111_11111110_00111100_01111110_01000000_10011010_11111111_11111111_11111111;
assign in[191] = 496'b00110000_00010001_01110111_00000101_11111111_01100101_00000010_11111111_10011111_01101011_11111000_11111111_00000100_01101011_11101010_00000100_01100111_11110001_11111111_11011110_01101110_01001000_01111101_10010001_11111111_11111111_11101111_00100001_01111101_01110000_11010100_11111111_10010000_01101110_01111011_01010010_01101110_00110001_11100010_00111111_01010101_10111110_11111111_11001101_01010000_01111000_01010001_00001000_00001000_00001000_00001000_01000000_01111101_10011000_00111010_01011000_01111110_01111110_01011000_11111111_11111111_11111111;
assign in[192] = 496'b11111111_11111111_11011100_01111011_00000110_11111111_11111111_11111111_10000010_01111101_00011111_11111111_11111111_11111111_11100010_01100110_01111101_11000110_11111111_11111111_11111111_00100110_01111101_01011001_11110011_11111111_11111111_11111101_01011100_01111101_10010011_11111111_11111111_11111111_10101011_01111101_01011111_11110101_11111111_11111111_10111100_01111001_01111101_10100011_11111111_11111111_11111111_00101011_01111101_01000001_11111010_11111111_11111111_11111111_01000010_01111100_11000010_11111111_11111111_00101110_11111111_11111111;
assign in[193] = 496'b01111011_10010110_11111111_11111111_11111111_01110110_01111010_11100111_11111111_11111111_11111111_11111111_00111010_01111011_11100111_11111111_11111111_11111111_11111111_10010111_01111010_11010011_11111111_11111111_11111111_11111111_11101000_01111011_10000010_11111111_11001110_10111001_11111111_11101000_01111010_01001001_01011100_01111011_01111010_11111111_11101000_01111011_01111100_01011101_00100001_01111011_11111111_11101000_01111010_01111011_01111010_01111011_01101100_11111111_11110010_01011101_01001010_00010111_10011011_11111111_11111111_11111111;
assign in[194] = 496'b11010011_01010011_01100100_00110011_00101001_11001110_01011111_01000011_11101001_11001100_01000110_11111111_01000100_01001001_11110100_11111111_11111101_10110110_11110101_01110100_00011110_11111111_11111111_11111111_11111111_11111111_00010010_01110111_10011101_11110001_11111111_11111111_11111111_11101110_00110010_01110001_01110010_01000000_11001000_11111111_11111111_11111111_11101001_10100011_00011011_01100100_11111111_11101011_10101000_10010000_10010001_00011011_00110101_11111000_01011111_01111011_01101111_01101111_01000000_11001110_11111111_11111111;
assign in[195] = 496'b01001101_01111100_01100101_01110100_01001010_10100011_01111101_10010100_11101001_01011111_01100001_11111111_00100111_01111101_11000000_00011111_01111100_10011011_11111111_10100101_01111101_01110010_01111100_00010100_11111111_11111111_11100010_01010000_01111101_01111101_00000001_11111111_10010110_01110010_01111101_00011001_00100000_01111100_10100101_01100001_01000010_11001000_11111111_11101000_01101001_01010100_01011000_11111000_11101111_10000110_01101111_01100101_11000010_01111100_01011100_01111101_01111000_00100000_11100010_10000001_11011010_11111111;
assign in[196] = 496'b11111111_10110011_01100001_10111011_11111111_11111111_11111111_10000011_01111011_10010101_11111111_11111111_11111111_11111111_10000011_01111011_11011000_11111111_11111111_11111111_11110110_01011100_01101110_11111000_11111111_11111111_11111111_10111101_01111101_00000000_11111111_11111111_11111111_11111111_00100100_01111100_10111100_11111111_11111111_11111111_11111111_00101010_01101111_11011100_11111111_11111111_11111111_11110111_01111011_00011101_11111111_11111111_11111111_11111111_11010010_01111011_10010000_11111111_11111111_01011011_11100011_11111111;
assign in[197] = 496'b11111111_11111111_11000100_01110110_11001110_11111111_11111111_11111111_00111111_01111100_11011110_11111111_11111111_11111111_11011110_01111110_00110000_11111111_11111111_11111111_11111111_10011011_01111101_10010010_11111111_11111111_11111111_11111111_01001011_01111000_11101110_11111111_11111111_11111111_11001101_01111100_00101101_11111111_11111111_11111111_11111111_10001111_01111110_10101100_11111111_11111111_11111111_11111111_01010010_01101111_11110001_11111111_11111111_11111111_11100000_01110100_00111100_11111111_11111111_01110110_10100110_11111111;
assign in[198] = 496'b11101101_01111100_00011001_11111111_11111111_11111111_11010110_01111110_10010010_11111111_11111111_11111111_11111111_10011101_01111110_11010111_11111111_11111111_11111111_11111111_00110010_01110001_11111111_11111111_11111111_11111111_11110011_01101001_00110001_11111111_11100001_00110101_11111111_11000010_01111110_10010100_10111100_01110001_01111100_11111111_00001010_01111110_01001110_01111110_01111110_10010111_11111111_00100010_01111110_01110111_01100100_11000101_11111111_11111111_11010111_10011010_11110000_11111100_11111111_11111111_11111111_11111111;
assign in[199] = 496'b11111111_11111111_11111111_11111111_11111000_01000111_10110101_11111111_11111111_11011001_01010000_11111111_11010001_01100100_11010011_10110101_01100100_01111000_11111111_11111111_10111010_01110101_01111110_01001110_10111100_11111111_11111111_10011101_00101010_11000101_11110101_11111111_11111111_11011010_01010010_11110110_11111111_11111111_11111111_11111111_00011110_10101100_11111111_11111111_11111111_11111111_11111111_01010011_11111101_11111111_11111111_11111111_11111111_11111111_01000101_11111111_11111110_11111111_11111111_00100000_01001110_10110001;
assign in[200] = 496'b00100001_01111000_01111110_01111110_01011100_10000110_01111111_00101101_11001110_00001011_01111110_11111111_10000110_01111110_00010010_11011001_01010101_01100101_11111111_11111010_01001011_01111110_01111100_01101010_11001111_11111111_11111110_00100001_01111110_01111110_00110100_11111111_11110110_00100111_01111101_00010111_01001001_01111100_11010111_01011110_01011110_11000101_11111111_10111010_01111110_10011101_00111000_01100110_10111000_11001100_01000011_01110111_11100010_11111000_00111100_01111110_01111110_01110110_10011100_10010000_10010011_11100000;
assign in[201] = 496'b01001111_01000000_10111101_11111110_11111111_01110000_10011101_00011000_01111101_10001011_11111111_00010111_01000111_00010111_01101100_01001000_01110010_11100101_11010101_00101001_00110010_10011101_11110001_01101011_10001011_11111111_11111111_11111111_11111111_11111111_00011010_00110100_11111111_11111111_11111111_11111111_11111111_00111000_00000110_11111111_11111111_11111111_11111111_10111101_01111101_11001000_11000111_11110101_11111111_11111111_00101111_01001101_11111100_11001000_00010001_11010000_00101000_01111010_10110101_01111110_01000010_10101111;
assign in[202] = 496'b01110011_00000110_00000110_01100100_11101000_01110001_11001001_11111111_11111111_00000011_10010000_11110110_01001111_11011111_11111111_11111111_00110100_10010000_11111111_11000001_01001000_11101101_10101001_01011000_11101000_11111111_11111111_10110000_01100111_01110000_10100111_11111111_11111111_11000000_00111101_00111100_00110001_01101011_10011000_10110010_01110001_10010111_11111111_11111111_11111011_00111001_01001100_10100011_11111111_11111111_11111111_11111111_11000010_10111100_01001101_10000100_10010011_00010011_01000011_10010000_10000001_10100111;
assign in[203] = 496'b01000110_00110101_10000010_01110000_10100010_01100111_11000011_11111111_11111111_00011110_00001100_10010100_00101111_11111111_11111111_11111111_01010101_10001000_11000000_01110010_11011101_11111111_11000101_01101011_11110100_11111111_10100010_01011001_00000101_01101000_10101010_11111111_11111111_11111111_11011000_01101000_01110100_00001001_11111001_11111111_11111111_00001010_00101010_11100100_00101111_01011101_11111111_11001100_01100100_11110110_11010101_00000010_01110001_11111111_10100000_01111110_01011110_01000111_10001110_10011110_10101000_11111111;
assign in[204] = 496'b11101000_00111001_01111100_01110011_01111110_11111111_00101111_01110100_10101000_11101101_01111110_11111111_11111111_01001000_01100010_11101100_00111001_01100011_11111111_11111111_10000001_01111110_01110010_01110010_11010010_11111111_11111111_10010001_01111101_01111110_10001000_11111111_11111111_10010100_01111010_01000100_01111001_01100111_11101111_00001101_01110110_10100000_11111111_10101011_01111101_10000011_01111110_10100111_11111111_11101100_10010110_01111110_10000111_00110011_01111011_01110010_01111001_01111100_00100111_10000001_10001100_11010100;
assign in[205] = 496'b10110001_00111001_01111000_01111101_01000111_00110110_01111101_01111011_01101000_01110101_01111101_10011101_01111101_01010010_11010011_11111111_11000010_01111101_00000001_01111101_10010000_11111111_10111100_01000001_01010001_10100111_01111101_01000111_00010000_01111010_01111101_10001100_11101111_01011110_01111101_01111101_01110110_10010000_11111111_11111111_00000111_01111101_01101000_10111011_11111000_11111111_11110100_01100010_01111101_00111100_01110101_00111110_11111111_10111010_01111101_01111101_01111101_01110100_10100100_01010010_10001001_11100110;
assign in[206] = 496'b11111111_11110111_01100001_11100001_11111111_11111111_11111111_11010000_01101000_11110100_11111111_11111111_11111111_11111111_00010110_10000010_11111111_11111111_11111111_11111111_11100010_01110001_11110101_11011101_11000110_11111111_11111111_00000001_00011010_10111001_01100101_00011010_11111111_11111110_01010001_00111000_01111001_10000011_11110100_11111111_11000010_01111110_01110011_10111011_11111111_11111111_11111111_00111001_01100001_11011110_11111111_11111111_11111111_11111111_00100110_11001001_11111111_11111111_11111111_11111111_11111111_11111111;
assign in[207] = 496'b11110000_01110110_11001110_11111111_11111111_11111111_11011101_01100101_11111111_11111111_11111111_11111111_11111111_10010011_00100111_11111111_11111111_11111111_11111111_11111111_00111000_10011011_11111111_11111111_11111111_11111111_11111000_01101000_11100101_11111111_11111111_10110011_11111111_11000011_01101000_11111111_11111111_11010100_01110011_11111111_10011100_00110110_11111110_10110101_01011110_01100110_11111100_01001011_01001100_01100010_01011000_10001001_11111000_11111011_10000001_10011110_11010000_11111101_11111111_11111111_11111111_11111111;
assign in[208] = 496'b01001010_01010010_00001000_01110001_00110010_10000011_01001111_11110010_11111111_11011100_10100011_11111111_01100001_11001011_11111111_11111111_11111111_11111111_11111111_01101000_11000101_11111111_11111111_11111111_11111111_11111111_00000010_01011101_10110110_11111111_11111111_11111111_11111111_11111111_10010110_01101100_01000010_10011000_11111111_11111111_11111111_11101101_00111001_01111101_00000100_11111111_11111111_11011100_01010110_00111100_11001001_11111111_11111111_11111111_00001011_01111101_00100001_01000110_00001101_10100111_10000001_10010000;
assign in[209] = 496'b10111101_01100111_11011001_11111111_11111111_01001101_00010110_00010010_10000100_11111111_11111111_11111111_11110111_00001111_01111010_01011011_11111111_11111111_11111111_11111111_11111110_00000110_01111000_11000000_11111111_11111111_11101011_11100101_00100100_00110100_01101000_11000101_11111111_10010000_01111101_00000011_11111111_10101001_01100101_11111111_00101011_00011000_11111101_11111111_11111100_01011011_11111111_10110110_01101010_10011010_00011011_01100001_01111101_11111111_11111010_00010110_01111010_01001111_00110010_11111111_11111111_11111111;
assign in[210] = 496'b11111000_01101111_01000010_11111111_11111111_11111111_10110001_01111110_10010100_11111111_11111111_11111111_11111111_00011001_01111110_11010011_11111111_11111111_11111111_11111000_01110010_01001111_11111111_11111111_11111000_11111111_10101111_01111110_00000110_11111111_11010110_01010010_11111111_00011011_01111110_11010110_10100100_01110011_01111110_11111111_01101011_01100111_00101101_01111110_01111101_10000111_11111111_01111101_01111110_01111110_01111110_00000010_11111111_11111111_01011111_00111000_00110001_10100101_11111111_11111111_11111111_11111111;
assign in[211] = 496'b10011011_01100100_01111101_01011010_11100010_00100111_00011000_11011101_11101100_00100111_00011110_11001110_01010000_11111011_11111111_11111111_10100000_01000110_10000010_10010110_11111111_11111111_11111111_10101010_00111100_00110001_10110100_11111111_11111111_11111111_00011101_00001001_00110001_11100111_11111111_11111111_11100111_01110011_11010010_00011101_10110100_11111111_11111111_00001001_00011110_11111111_11001001_10001011_11111111_11000100_01101110_11100111_11111111_11111111_00011101_00110110_01010101_10101010_11111111_01101001_10000110_11111111;
assign in[212] = 496'b01010001_10100111_11001011_11111111_11111111_01011000_11101110_11111111_11111111_11111111_11111111_00011000_00001010_11111111_11111111_11111111_11111111_11111111_10111011_01101010_01000111_10101000_11111110_11111111_11111111_11111111_11101010_10001110_01111010_10110111_11111111_11111111_11111111_11111111_11111101_01011111_11010001_11111111_11111111_11111111_11111111_10101100_01010111_11111100_11111111_11111111_11111111_11111111_10110011_01110111_11010001_11111111_11111111_11111111_11111111_11111111_00000101_01110100_01001110_11111111_11111111_11111111;
assign in[213] = 496'b01010001_11100010_11111111_11111111_11111111_11111111_00110100_11000100_11111111_11111111_11111111_11111111_11111111_00001010_10001110_11111111_11111111_11111111_11111111_11111111_10001011_10001011_11111111_11111111_11111111_11111111_11111111_10001011_01011000_00011111_00101110_11001010_11111111_11111111_00101011_10111011_11111111_11100111_00100111_11111111_11110111_01101011_11100101_11111111_10110001_10001001_11111111_11101010_01111110_11100101_11010110_01010101_11100101_11111111_11110110_10001100_01001100_00110111_11100010_11111111_11111111_11111111;
assign in[214] = 496'b11111111_11000100_01110111_00111110_11111111_11111111_11111111_00011101_01111101_00010010_11111111_11111111_11111111_11111111_01010000_01111101_10100110_11111111_11111111_11111111_11010011_01111000_01111101_11101010_11111111_11111111_11110011_01011101_01111101_01111101_10101100_11111111_11111111_11101011_01111101_01111101_01110111_11010001_11111111_11111111_11100000_01111101_01111101_01001011_11111111_11111111_11111111_10010001_01111101_01111101_10100000_11111111_11111111_11111111_00100000_01111101_01110110_11101011_11111111_10001011_10111111_11111111;
assign in[215] = 496'b11111111_11010111_10100011_10000001_10110111_11101001_00010001_01110110_01111101_01111110_01111100_10100111_01101010_01111110_01111110_01010111_10010010_01111110_01111101_00111101_00101001_01111100_10111101_00001010_01111000_00111000_10011000_01110100_10011000_11110101_01100100_01010010_01110110_01100100_00011111_11111111_10011000_01111110_01010111_11110001_11111101_11111111_11111111_00110000_01111110_01100100_11111111_11111111_11111111_11101011_01101010_01111100_10101100_11111111_11111111_11111111_00001011_01111110_10001100_11110011_01110010_00110111;
assign in[216] = 496'b11111111_11111111_11111111_11111111_11111111_00010111_11111111_11111111_11111111_11111111_11111111_01010011_00010111_11111111_11110111_10111011_10001010_10011000_01100101_10000011_10011101_01011100_01100011_00011011_00111101_01111110_01011001_01000111_11000110_11111011_11111111_10011001_01110101_10010100_11111111_11111111_11111111_11111111_00100111_10001011_11111111_11111111_11111111_11111111_10101100_01110000_11111111_11111111_11111111_11111111_11101101_01100100_00000001_11111111_11111111_11111111_11111111_00101001_00111101_11111111_11111011_01010101;
assign in[217] = 496'b10111011_01101001_10100110_00100010_10101010_11000010_01110001_10101011_11100111_01011100_10101111_11111111_00000101_00001001_11111111_10000011_00110001_11111101_11111111_00000101_00111110_10011011_01010000_11011010_11111111_11111111_11100010_00110111_01111101_01100010_11001001_11111111_11111111_11111111_00001010_10101101_00101100_01110100_11001100_11111111_10011101_10110101_11111111_10011000_01111101_10111000_11000100_00010100_11110010_10011101_01001111_10000010_11111111_10101110_01101111_01010110_01011011_10010101_11111111_10000010_11110100_11111111;
assign in[218] = 496'b11111111_11111110_10011101_11111111_11111111_11111111_11111111_11010010_01110111_11110100_11111111_11111111_11111111_11111111_00011011_00111000_11111111_11111111_10001011_10001001_00000010_01111001_00110010_10011010_00100010_01110100_01111110_01111110_01111110_01111110_01111110_01111110_11111001_11010001_01110001_00001101_11001111_00011111_01110110_11111111_10010000_01101111_11110100_11111111_01000001_00010100_11111001_01011011_10000010_11111111_11111111_11101010_11111001_11101100_00001000_11110110_11111111_11111111_11111111_11111111_11111111_11111111;
assign in[219] = 496'b11110101_11111111_11111111_11111111_11110011_01111110_01111000_00110110_11110001_11110101_01001011_01101111_00100110_01101000_01111110_01000011_00001111_01111110_11010111_11111111_11111010_01000010_01111110_01111110_00101110_11111111_11111111_11111111_11011011_01111001_01100000_11101111_11111111_11111111_11111111_00011001_01111110_10110111_11111011_11111111_11111111_10111001_01110100_01001110_10001111_01011001_11111111_11111111_01000000_01111110_01111110_01111110_01011011_11111111_11101111_01111001_01111110_01010111_10111000_10111110_11001110_11111010;
assign in[220] = 496'b11111111_11000011_00101101_01111001_01101011_11111101_00001101_01111000_00010111_11010000_11010011_11111110_00100101_01001111_11010011_11111111_11111111_11010011_00000000_01011000_11101101_11111111_11111111_11111111_10000001_01011010_11011101_11111111_11111111_11111111_11111101_01001010_00000000_11111111_11111111_11111111_11111111_10101011_01010011_11001101_11111111_11111111_11111111_11011110_01100001_11000011_11001101_11111111_10110010_00100100_01111000_00000100_11111111_00001101_11011111_10011011_01111100_01000111_11111101_00110101_00000001_11110011;
assign in[221] = 496'b11111111_10011111_01011000_11111111_11111111_11111111_11111111_01000011_10001110_11111111_11111111_11111111_11111111_11011100_01111010_11010100_11111111_11111111_11111111_11111111_10100010_01010010_11111111_11111111_11111111_11111111_11111111_01000110_00000100_00100100_00101000_11111111_11111111_11010110_01100010_01101000_10100011_00101110_10100010_11111010_00011001_01001110_11011001_11111111_00001000_00000010_10101011_01110011_11010011_11101110_00101011_01001010_11100101_11111011_10111100_10101010_01011100_00000110_11101111_11111111_11111111_11111111;
assign in[222] = 496'b00100100_01000111_01011010_01100001_10100010_01011101_10010110_11110011_11111111_11100101_00001010_01100111_11010010_11111111_11111111_11111111_11111111_11111111_10010010_01011010_10111100_11111110_11111111_11111111_11111111_11111111_10101010_01001000_01010000_10000100_10100101_11111011_11111111_11111111_11111111_00000001_01111101_00111101_11110000_11111111_11111111_10101011_01001000_11010001_11111111_11111111_11111111_11110100_01100110_11100100_11111111_11011010_00111001_11111111_11000001_01001101_11110001_11000011_01011100_00111101_01111111_01011111;
assign in[223] = 496'b00010000_01111111_01100000_00010000_11111111_11111111_01111111_11000000_11111111_10110000_11111111_11111111_11111111_01100000_10110000_11111111_11111111_11111111_11111111_11111111_00000000_01100000_11110000_11111111_11111111_11111111_11111111_11110000_01100000_00101111_11111111_11111111_11111111_11111111_11111111_00010000_01111111_10010001_11111111_11111111_11111111_10010001_01101111_00100000_11100000_11111111_11111111_11111111_00000000_01000000_11110000_11111111_11111111_11111111_11111111_11110000_01000000_01101111_00100000_11111111_11111111_11000000;
assign in[224] = 496'b11111111_11101011_10011110_00011010_10100101_11111111_11000011_01101010_00001000_10001110_00110111_11111111_11111111_00110000_10000010_11111111_11111111_11010110_11111111_11111111_00001110_00010010_11111110_11111111_11011001_11111111_11111111_11011101_01100101_10110011_11111111_11111111_11111111_11111111_11111111_10100001_01001101_11111111_11111111_11111111_11111111_11111111_11111000_01011100_11011000_11111111_11000100_11010111_00001110_10000010_01101000_10000111_11111111_00011011_00011011_00000010_00011011_10101010_11111110_11111111_11111111_11111111;
assign in[225] = 496'b10111110_00100110_01000011_01011001_10111111_11001000_01101111_10010100_11011101_11100101_11111111_11111111_10100011_01000010_11110101_11111110_11111111_11111111_11111111_11101100_00111110_01101111_01011001_11101101_11111111_11111111_11111111_11111111_11011010_01010001_11101001_11111111_11111111_11111111_11111111_11111111_00010101_10110000_11111111_11111111_11111111_11111111_11111111_00010101_10100101_11111111_11111111_11111111_11111111_11111111_00010101_10010011_11111111_11111000_11100100_11111111_11100000_01001000_10110111_00110111_01110000_00001101;
assign in[226] = 496'b11000110_00100111_01111010_01111110_01011111_11001110_01111000_01100110_00000001_00100100_01111110_11111111_10010000_01111110_10011100_11010011_01110010_00101100_11111111_11010111_01110011_01101100_01101001_01001000_11110000_11111111_11111111_10000011_01111110_01111110_11010001_11111111_11111111_11000001_01101000_01100110_01111101_00101101_11111111_10011101_01110111_01000010_11110001_00010101_01111100_11100111_01110110_10001000_11111001_11110011_00101110_01111011_11100100_01101010_10100011_00010101_01100110_01101100_10101011_01001100_10010000_11101011;
assign in[227] = 496'b11111111_11001101_10001101_11011101_11111100_11111111_11010100_01100100_01111110_01111101_01001101_11111111_00000001_01111000_01111101_01111101_01101111_01111110_10001001_01111101_00110111_01011111_01110011_00100111_01111110_01110101_00100100_10100000_01111101_00000101_01100010_01011010_01111101_00010000_01111101_00111111_10101001_01111101_10000001_01111101_01111010_00000100_11111111_01011001_01101101_11100001_10100111_11101011_11111111_11010010_01111101_00100111_11111111_11111111_11111111_11111111_10000011_01111101_10111011_11111111_00010111_01111101;
assign in[228] = 496'b11010101_00100001_01001000_01110101_00011001_10101111_01110000_10000100_11011101_00100000_00101110_11111111_01001011_11010110_11111111_00000011_01011011_11101010_11111111_11111111_11111111_10011011_01010010_11100100_11111111_11111111_11111111_10111011_01101001_11010100_11111111_11111111_11111111_11111100_01010011_10000111_11111111_11111111_11111111_11111111_11000101_01110110_11110111_11111111_11111111_11111111_11111111_11000101_01001000_11111111_11111111_11111111_11111111_11111111_11010100_01101111_10111011_10110010_00011111_10001100_01110111_01010100;
assign in[229] = 496'b11111111_11111111_11111111_11111111_11111111_11001100_11111111_11111111_11111111_11111111_11111111_11101010_00111100_10001000_11001010_11111010_11111111_11111111_11111111_11111010_10111011_00000010_01101001_11100100_11111111_11111111_11111111_11111111_10000111_00011000_11111111_11111111_11111111_11111111_11001001_01000000_11111010_11111111_11111111_11111111_11111111_00111001_11010100_11111111_11111111_11111111_11111111_11111111_10110010_00110101_00111001_00100100_00001001_11111111_11111111_11111111_11111111_11111100_11100110_11111111_11111111_11111111;
assign in[230] = 496'b01100101_11001101_11111111_11111111_11111111_01100100_11010010_11111111_11111111_11111111_11111111_01000001_10001011_11111111_11111111_11111111_11111111_11111111_00011101_11000011_11111111_11111111_11111111_11111111_11111111_00011000_11000100_10101010_10000010_10000010_10000010_10101010_10000001_01111101_00110111_10000001_10000001_00010011_01000110_11110110_01000110_10010110_11111111_11111111_11101100_00001001_11111111_11100010_01010000_00010011_10001100_01001011_00011110_11111111_11111111_11100111_10001011_10010110_11100010_11111111_11111111_11111111;
assign in[231] = 496'b01101100_00110000_00000000_11110111_11111111_00100111_00001111_11111111_11111111_11111111_11111111_11111111_01001001_10001111_11001101_10101110_11110000_11111111_11111111_10111111_00110100_01000001_01100000_01100110_10110111_11111111_11111111_11111111_11111111_11111111_10010101_00110111_11111111_11111111_11111111_11111111_11111111_10011011_00111000_11111111_11111111_11111111_11111111_11111110_01000011_10011010_11111111_11111111_11110110_11011101_10100100_01111101_11010110_00001100_01010010_01110001_01101100_00101011_10000101_11001001_11110111_11111111;
assign in[232] = 496'b01010000_01101000_11110101_11111111_11111111_11011000_01111110_00001111_11111111_11111111_11111111_11111111_00010001_01111110_11011111_11111111_11111111_11111111_11111111_01000010_01111001_11111100_11111111_11111111_11111111_11100001_01111110_00100111_11111111_11111111_11000110_01000110_11001101_01111110_10001010_11101011_00011110_01110100_01111110_10101011_01111110_01000111_01110000_01111110_01110101_10001011_10100000_01111110_01111110_01111110_01011110_11011010_11111111_11101111_10000101_10110000_10100001_11111100_11111111_11111111_11111111_11111111;
assign in[233] = 496'b11110100_10011011_00101111_00000101_11010000_11100111_01100101_01111101_01011101_01111110_01110000_11111111_10001100_01110001_11011101_11111101_00101000_10101110_11111111_10011100_01111101_00010110_10000010_00101100_01011001_11111111_11111001_10001011_01001101_01010110_01011010_01111101_11111111_11111111_11111111_11111111_11111111_01001000_00111110_11111111_11100111_10110010_10001000_01001001_01101111_11011010_01010111_01111100_01111110_01111000_00110111_10110000_11111111_00001110_10101110_11001101_11110010_11111111_11111111_11111111_11111111_11111111;
assign in[234] = 496'b11111010_00010111_01111001_01111101_01000111_11111111_00011010_01111101_00010100_01110101_01100101_11111111_11101001_01111010_00000011_10101111_01111101_00000011_11111111_11101110_01111001_11001011_01101000_01101001_11111110_11111111_11111111_00111010_01101001_01111100_10101100_11111111_11111111_11110101_00111110_01111101_10010110_11111111_11111111_11011111_01000001_01100100_00100101_00110111_11111110_11111111_10101100_10110010_11100101_10100001_01111101_10101011_11111111_00010000_00101110_01011100_01111101_01110111_11001000_10000001_10000001_11001110;
assign in[235] = 496'b11010001_01111010_01001000_11111111_11111111_11111111_10001111_01111110_10100100_11111111_11111111_11111111_11111101_01011101_01011111_11111100_11111111_11111111_11111111_11010101_01110111_00101000_11111111_11111111_11111111_11111111_00001011_01111110_10110100_11111111_11111100_10100110_11111110_01100000_01101101_11101000_11011001_01000001_01111101_11101101_01111110_00111011_00000010_01110000_01111110_00101011_11101101_01111101_01111110_01111101_01100101_11000111_11111101_11101101_01111110_01101011_00111000_11100011_11111111_11111111_11111111_11111111;
assign in[236] = 496'b00011111_01110100_01110100_00111110_00111110_00101011_01101011_10010010_11110010_11111111_11111111_11111111_01001000_10010111_11111111_11111111_11111111_11111111_11111111_00110000_01100101_10000111_11101001_11111111_11111111_11111111_11110000_00001110_01110011_01111000_00111100_10101001_11111111_11111111_11111111_11100101_10001101_01111101_01111100_11111111_11111111_11111111_11111111_10110110_01111101_00100011_11111111_11111111_11111111_11111111_11111010_00110100_11011111_00111110_00111101_00111101_00111110_00111010_11101111_10010011_10110110_10111001;
assign in[237] = 496'b11111111_11111111_00100010_01111110_11010010_11111111_11111111_11100111_01111001_01010101_11111011_11111111_11111111_11111111_10010001_01111101_10000110_11111111_11111111_11111111_11111111_01000110_01111101_11111011_11111111_11111111_11111111_11011000_01111000_01010101_11111111_11111111_11111111_11111111_10011011_01111101_10000001_11111111_11111111_11111111_11111111_00101100_01111101_10111001_11111111_11111111_11111111_11111111_01101110_01101110_11111111_11111111_11111111_11111111_11111111_01111101_01001011_11111111_11111111_10001011_10111001_11111111;
assign in[238] = 496'b11111111_11111111_11101111_10110101_10011000_11111111_10101100_00100010_01111010_01101011_01101101_11111101_00100001_01111100_00111101_11000000_11111000_11101100_00101111_01101111_10100111_11111111_11111111_11111111_11111111_01101000_11001011_11111111_11111111_11111111_11111010_00001000_00110000_11111111_11111111_10001100_10110000_00111111_01111101_01010001_10011000_11010100_00100011_01111101_01011100_10100001_01110001_01111101_01111101_01111101_00100111_11110011_11111111_11101000_10101101_10010111_11000110_11111111_11111111_11111111_11111111_11111111;
assign in[239] = 496'b11111111_11000000_01110001_11001001_11111111_11111111_11111111_01000101_01011111_11110001_11111111_11111111_11111111_10111100_01111111_10010010_11111111_11111111_10001011_00010111_01010010_01111110_00011011_00010111_10001011_01100100_01001111_01111110_01001000_00101110_01100000_01111110_11111111_10011110_01111101_11011110_11111111_11011000_01111110_11111111_00110001_01000000_11111111_11111111_01001000_01001010_11101010_01110111_10001111_11111111_11111111_00110010_11101010_10100110_01110011_11110001_11111111_11111111_11100111_11111111_11111111_11111111;
assign in[240] = 496'b11111111_11111111_11110011_10010111_00100111_11111111_11111111_10011010_01011100_01001111_00011110_11111111_11101100_00101110_01010111_11000111_11111111_11111111_11100011_01010011_00011001_11110100_11111111_11111111_11110001_01011101_00001000_11111111_11111111_11111111_11111101_00011001_01101111_11111001_11100110_11111101_11111101_00011000_01110000_10001111_11111111_11011101_00101001_01001101_01101001_11001111_01000110_00010001_01100101_01111011_00110101_11101100_11111111_01010111_01011011_00101000_11010010_11111111_11111111_11111111_11111111_11111111;
assign in[241] = 496'b11111101_10100010_01010101_01111101_01011100_11111010_10001010_01111101_01111101_01001101_01111101_10000101_01001110_01111101_01111101_01111101_01101000_01111101_10111011_01111101_01111101_01111101_01111101_01111101_00100111_10000111_01111101_10011010_11101101_11101101_11101101_11111011_01101101_01011011_11110111_11111111_11111111_11111111_11111111_01111101_01010011_11111111_11111111_11111111_11111111_11111111_01111101_01010011_11111111_11111111_11110101_00000110_11000010_00000100_01110111_00001000_11100101_00110010_01111101_01111110_01111110_01111110;
assign in[242] = 496'b11110111_10101110_10000010_10101001_11111110_00001101_01110110_01100110_01111100_01111101_00100010_00101000_01010100_11000111_11111001_10110111_01111000_01111101_01111000_10101010_11111100_11011010_00011011_01111101_01111100_01001101_01111001_01010011_01111101_01111100_01111101_01100100_11100001_00011001_10001100_11001010_00010010_01111110_10000010_11111111_11111111_11111111_10001111_01111100_00010111_11111111_11111111_11111111_10100010_01110111_00100100_11110100_11111111_11111111_10011110_01110101_10001011_11111111_11111111_10001100_11111111_11111111;
assign in[243] = 496'b11111111_11111111_01001001_01110111_11010001_11111111_11111111_10100110_01111101_00000100_11111111_11111111_11111111_11110100_01100100_01011000_11111010_11111111_11111111_11111111_10101111_01111100_10110010_11111111_11111111_11111111_11111111_01001111_01000101_11110111_11111111_11111111_11111111_10110010_01110111_10110101_11111111_11111111_11111111_11110100_01001011_00101100_11111111_11111111_11111111_11111111_11001000_01111001_11011010_11011110_10010011_00010010_10011111_11010100_01111010_01100010_01000101_01000101_01000101_11111111_11111111_11111111;
assign in[244] = 496'b01111100_01111101_00111011_11111111_11111111_01111110_01000111_00111111_01011111_11111000_11111111_11001100_01111101_11010011_00001100_01101010_11110000_11111111_11110111_01100110_01001110_01100100_00010100_11111100_11111010_11111111_11010101_01110110_01111110_01100100_00110100_01100001_11111111_10110000_01111001_00100111_01011010_01100101_01111101_11111111_00111001_00111010_11111111_10110111_01111101_01001011_11111111_10000010_01111100_00101111_01000010_01111010_10000011_11111111_11100011_01000010_01111101_01111010_00000001_11111010_10100000_11010001;
assign in[245] = 496'b11111111_11111111_11111111_11111111_11111111_11111111_11111101_00010111_01010101_01001010_00010011_11111111_11111111_11000011_01010011_11010010_11101000_10011111_11111111_11111111_10101111_01000111_11111100_11111111_11010001_11111111_11111111_11111001_01011100_10000011_11111001_11111111_11111111_11111111_11111111_10101000_01111110_01011101_11111011_00000101_00001001_00010000_01111010_00100011_11100101_11111111_00000101_10011010_00001000_00000010_11011101_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111;
assign in[246] = 496'b11111111_10100101_00110110_11111111_11111111_11111111_11111111_01010011_10100010_11111111_11111111_11111111_11111111_11010100_01110111_11101011_11111111_11111111_11111111_11111111_00010011_00101000_11111101_11100001_11111101_11111111_11101001_01111101_00000100_01001000_01101110_10111001_11111111_00000010_01111110_00001110_11101101_01011001_11001110_11101000_01110101_00000011_11111111_10011000_01010100_11111100_11111111_00111110_10010111_00011111_01001001_11011101_11111111_11111111_11011101_10000001_10110101_11111100_11111111_11111111_11111111_11111111;
assign in[247] = 496'b00000010_11111111_11111111_11111111_11111111_00110100_00010011_11111111_11111111_11111111_11111111_11111111_00110011_01101101_00101101_10010100_11111010_11111111_11111111_01101111_00011111_10001110_01010000_01001111_11100110_11011110_01111011_11010111_11111111_11101110_01010000_00111110_10010001_01101000_11110101_11111111_11111111_10001000_01101111_00011110_10101010_11111111_11111111_11111111_10011001_01101111_11001011_11110010_11111111_11111111_11111111_10001011_01001011_11111111_11111111_11111111_11111111_11111111_11001011_11111111_11111111_11111111;
assign in[248] = 496'b11111111_11111111_11110101_10101010_11111100_10010011_11111111_11111100_00100000_01011111_11100101_11111111_00110110_00011101_00110101_01100000_00011111_11111111_11111111_11111110_00000111_00100001_11001101_11111111_11111111_11111111_11111111_00101100_11101110_11111111_11111111_11111111_11111111_11000111_00010000_11111111_11111111_11111111_11111111_11111111_10011001_10100001_11111111_11111111_11111111_11111111_11111111_11100100_00100111_11111100_11111111_11111111_11111111_11111111_11111111_10010110_10000101_11111111_11111111_11111111_10100010_10000001;
assign in[249] = 496'b11111111_11111111_10110100_01111101_00110101_11111111_11111111_11101010_01101100_01111101_10100011_11111111_11111111_11111111_10010001_01111101_00100011_11111111_11111111_11111111_11111111_01011111_01111011_10110001_11111111_11111111_11111111_11101010_01110101_01010101_11111111_11111111_11111111_11111111_10100001_01111101_00101000_11111111_11111111_11111111_11111111_00110001_01110101_11010111_11111111_11111111_11111111_11011101_01111100_01010001_11111111_11111111_11111111_11111111_00001000_01111001_11010010_11111111_11111111_10101000_11111111_11111111;
assign in[250] = 496'b10111001_01101001_00111100_00110010_01111001_11001110_01101001_10011111_11111111_11100010_01111001_11111111_00011000_00001110_11111111_11101100_01010000_00110010_11111111_00010011_00000100_11111011_01000110_01010000_11101100_11111111_11011101_01111000_01001011_01000110_11101100_11111111_11111111_11110001_01101001_01111101_11100111_11111111_11111111_11111111_00010011_01101001_01111000_10100000_11001001_11111111_11011101_01111000_11001000_10010101_01101110_01000001_11100010_11011101_01111000_00010011_00000100_01101001_01010000_10000001_10000001_10001011;
assign in[251] = 496'b01001001_11111111_11111111_11111111_11111111_11111111_01010000_11111111_11111111_11111111_11111111_11111111_11101011_01000000_11111111_11111111_11111111_11111111_11111111_11100010_01101010_00111011_01001011_01011000_11110010_11111111_11100010_00011011_11111111_11111111_00010110_11100010_11111111_10110100_10010101_11111111_11111111_00110010_11111111_11111111_10010010_10101110_11111111_11110101_01000110_11111111_11111111_00001110_10111000_11111111_10111111_00001010_11111111_11111111_00010110_11110111_11111111_10010111_10100000_11111111_11111111_11001110;
assign in[252] = 496'b11111111_11100111_01000011_01101101_00110110_11111111_11111111_00101000_01110001_10010101_01111110_11111111_11111111_11111111_00110100_01000001_10110000_01111101_11111111_11111111_11111111_00011011_01101011_01101111_00010001_11111111_11111111_11101001_01011000_01110011_11001001_11111111_11111111_11100111_01010100_01101101_01111000_11100111_11111111_11010000_01101101_00011111_11100011_01111101_10111011_11111111_01101001_00010001_11111100_11011111_01111110_11010100_11111111_00100100_11111100_10011110_01010000_00101100_11111111_00010001_00000000_11111100;
assign in[253] = 496'b11011110_01000001_01110011_01001001_00000101_11100011_01101000_00111011_10010011_00001011_01010101_11111111_10000111_01100101_11111110_11111111_11111111_11001011_11111111_00101000_00011100_11111111_11111111_11111111_11111111_11111111_00001110_00011110_11111111_11111111_11111111_11111111_11111111_10100101_01110110_00100101_11011001_11111111_11111111_11111111_11110110_01100011_01010111_11010101_11111111_11111111_11111111_11111111_01010110_10000100_11111111_11111111_11111111_11111111_11111001_01101110_00001110_00000001_01010100_10101000_01101010_01101010;
assign in[254] = 496'b11101100_10001111_10000001_11010100_11111111_11100010_01000110_10000011_01010001_01011010_11111000_11111111_00111010_10111000_11111111_11101110_01111001_11101101_11111111_01011110_01001000_10100000_10100101_01111001_11011011_11111111_10101000_00101100_01011011_01100000_01011010_11111110_11111111_11111111_11111111_11111110_10010111_10000011_11111111_11111111_11111111_11111111_11101110_01010000_11100100_11111111_11111111_11111111_11111111_00010010_00100010_11111111_11111111_11111111_11111110_10100011_01100110_11110001_11111111_01101111_10111111_11111111;
assign in[255] = 496'b01010100_11111010_11111111_11111111_11111111_10011100_01111011_01010111_00101000_01100110_00111101_11111111_11111100_01000010_01111100_01111101_01111100_01111100_11111111_10100111_01111011_10110000_11011010_10001111_10000111_11111111_01100100_00110000_11111111_11111111_11111111_11111111_10111100_01111100_11001101_11111111_11111111_11111111_11111111_10011000_01110001_11110001_11111111_11111111_11111111_11111111_10011000_01111100_11011011_11111111_11111111_11111111_11111111_11010000_01111011_00010010_10110100_10110011_10000111_01101011_01111101_01111010;
assign in[256] = 496'b00100011_11111111_11111111_11111111_11111111_00110100_00100000_11111111_11111111_11111111_11111111_11100101_01110100_10011100_11111111_11111111_11111111_11111111_10011101_01111101_11010000_11111111_11011111_00110010_00111111_10010000_01111100_00001001_00001100_01111101_01100101_01001110_10011010_01111100_01111100_01101111_10001111_11100101_11011111_11111011_00010000_01110010_11010101_11111111_11111111_10101000_11111111_11111011_01001000_01010010_10110001_00011100_01101111_11111111_11111111_11101001_01000001_01111110_01110001_11111111_11111111_11111111;
assign in[257] = 496'b11101100_10010010_10010111_11101000_11111111_11010001_01110110_00110010_00111010_01011011_11111111_11011001_01011011_10110010_11111111_11111101_01001111_10110001_10001101_00001011_11111111_11111111_11111111_00110010_10001101_11010110_01100010_00010001_00010001_01001111_01111010_10111111_11111111_11010011_10001111_10011110_10010011_01111011_11111110_11111111_11111111_11111111_11111100_00111101_00000000_11111111_11111111_11111111_11111111_00000001_01100000_11100001_11111111_11111111_11111111_10100110_01101111_11010001_11111111_01011011_11000111_11111111;
assign in[258] = 496'b11111111_10111110_01101001_01111101_01011111_11111111_11100111_01101001_00110010_10110100_01101001_11111111_11111111_11010011_01110100_11010111_00011000_01101110_11111111_11111111_11010011_01111000_00111011_01111000_11000011_11111111_11111111_10111110_01111101_00111100_11101100_11111111_11111111_11000100_01100100_01001011_01011111_11110001_11111111_11010011_01101001_01001100_11101100_01011111_00010011_11111111_01000001_01010110_11110001_11100111_00101100_00110010_11111111_01111001_10010110_01010000_01101110_01101110_11001110_11111111_11010010_11110001;
assign in[259] = 496'b11111111_01010011_00111011_11111111_11111111_11111111_11111111_01001001_01010000_11111111_11111111_11111111_11111111_11111111_01001001_01110110_11111111_11111111_11111111_11111111_11111111_01001001_01110110_11111111_11111111_11111111_11111111_11111111_01110101_01010100_11111111_11111111_11111111_11111111_11111011_01111011_00011100_11111111_11111111_11111111_11111111_10011101_01111101_11010011_11111111_11111111_11111111_11111111_00101101_00110001_11111111_11111111_11111111_11111111_11111111_01010111_00001111_11111111_11111111_01101101_11101000_11111111;
assign in[260] = 496'b01110011_00011000_11111111_11111111_11111111_11111111_00101100_00011000_11111111_11111111_11111111_11111111_11111111_01011111_10000110_11111111_11111111_11111111_11111111_11001101_01111101_11100010_11111111_11111111_11111111_11111111_11000011_01111101_11111111_11111111_11111111_11111111_11111111_00000100_00110110_11111111_11111111_11111111_11111111_11111111_01000001_10011011_11111111_11111111_11111111_11111111_11111111_00101100_01011111_01011111_01111101_01111101_01111101_11111111_00011000_00000100_11110110_11111111_11111111_11111111_11111111_11111111;
assign in[261] = 496'b11111111_11100010_00100011_01110011_01111101_11111111_10101100_01100010_01011110_00010011_00111101_11111111_10001100_01111100_00100011_11110011_11111111_10110011_11000011_01110100_00110101_11111110_11111111_11111111_00010011_00100110_01100100_11101101_11111111_11111111_11101100_01101101_01111011_10011001_11111111_11111111_11111110_00111001_01011111_01111101_10110010_11111111_11111110_00001111_01111100_00000001_01110111_10011011_11110100_00100110_01111101_00011110_11111111_01100011_01110100_00011111_01111101_01011001_11111000_01111001_01010101_10001000;
assign in[262] = 496'b11111111_10000100_01111101_10011101_11111111_11111111_11111111_00111011_01100000_11111101_11111111_11111111_11111111_10110011_01111101_10010000_11111111_11111111_11111111_11111111_00101100_01010110_11110100_11111111_11111111_11111111_11101101_01110001_10000100_11111111_11111111_11111111_11111111_10101011_01111101_11001110_11111111_11111111_11111111_11111111_10001011_01101011_11111001_11111111_11101000_11110110_11111111_10001011_01110110_00010000_01011110_01111000_01101111_11111111_10101101_01111001_00101111_10000101_00000000_11111111_11111111_11111111;
assign in[263] = 496'b11111111_00001111_00100111_11111111_11111111_11111111_11101001_01110000_11001100_11111111_11111111_11111111_11111111_00001000_00100111_11111111_11111111_11111111_11111111_11110111_01100100_11001011_11111111_11111111_11111111_11111111_10111100_01010011_10100100_00110100_01000011_10011110_11111111_10001001_01101000_10001011_11011101_10100000_01001010_11111111_00011101_11001110_11111111_11011110_01010110_10101110_10001100_11110111_11111010_10011111_01101001_10010101_11111111_10011110_01001001_00111100_00011111_11010100_11111111_11111111_11111111_11111111;
assign in[264] = 496'b00111010_01100101_00110010_11001100_11111111_11111111_00111010_01101010_00000111_01011101_00101011_11111111_11111111_00001011_01100011_11111111_11110110_00001011_11111111_11111111_10010001_01110110_11111111_11111111_11011110_11111111_11111111_11011010_01111100_11011110_11111111_11111111_11111111_11111111_11110011_01110000_10101101_11111111_11111111_11111111_11111111_11111111_00111110_10000110_11111111_11111111_11111111_11100101_11111111_00101010_00100110_11111111_11111111_11111110_01110100_01000000_01100100_00110001_11111111_00100000_01101100_00011011;
assign in[265] = 496'b11111111_11111111_11111111_11111111_11111111_00001111_01100010_01111101_01100011_00000101_11101111_00000001_00111010_10111011_11010110_10111100_01001000_00101111_01001011_10010001_11001011_11110000_10100011_00011001_01011101_10110100_01010011_01110010_01010111_00110111_01101100_00110010_11111111_11111111_11111111_11111111_11111111_01000110_10110000_11111111_11111111_11111111_11111111_11000100_01110111_11100110_11111111_11111111_11111111_11110111_01000000_10000011_11111111_11111111_11111111_11111111_10100000_01100110_11100100_11010011_01101001_10100111;
assign in[266] = 496'b10000010_11010110_11111111_11111111_11111111_10101001_01010100_01111100_00000010_11111101_11111111_10110110_11111111_11010010_10000011_01111001_00101101_11111111_10000100_11111111_11111111_11111111_10100001_01110000_11110100_01000011_10010100_11011000_11000010_00111000_01111101_10010001_11101101_00100100_01101001_01100000_10000110_00001110_00011001_11111111_11111111_11111111_11111111_11111111_10000010_00111110_11111111_11111111_11111111_11111111_11111111_00001010_00111110_11111111_11111111_11111111_11111111_11111011_01010110_01010111_00001001_01001110;
assign in[267] = 496'b01111101_01110101_00001110_11111000_11111111_01001110_10001010_00010110_01111001_01011011_11000101_01111100_10101010_11111111_11111111_11000111_01101101_01011010_01110000_11111100_11111111_11111111_11111111_10110010_01111100_01111101_10111011_11111111_11111111_11111111_11111111_01101110_01100000_00101111_11111010_11111111_11111111_11011000_01111100_11011100_01100000_00011000_11111111_11111111_10010000_01111101_11111111_00000010_10010101_11111111_10111110_01100011_01011010_11111111_00000100_01010001_00111011_01111001_01100110_00101101_01100111_00011101;
assign in[268] = 496'b11011011_00111001_11110111_11111111_11111111_11111111_11110111_01011110_11101010_11111111_11111111_11111111_11111111_11101010_01111101_11010100_11111111_11111111_11111111_11111111_11101010_01111101_11101010_11111111_11111111_11111111_11111111_11101010_01111110_11101010_11111111_11111111_11111111_11111111_11101010_01111101_11101010_11111111_11111111_11111111_11111111_11101010_01111101_11101010_11111111_11111111_11111111_11111111_11101010_01111101_11101010_11111111_11111111_11111111_11111111_11101110_01110100_11101010_11111111_11111111_00110011_11101010;
assign in[269] = 496'b00101001_01001001_00001001_01011100_00001100_00001110_01010110_11110000_11111111_11011010_01101101_11110101_01011101_11100001_11111111_11111111_11111111_00110011_11100101_01011111_11111111_11111111_11111111_11111111_00110011_11010110_00101010_11111111_11111111_11111111_11111111_00111000_10101100_01011110_11110000_11111111_11111111_11111000_01101100_10101100_01011111_00000001_11111111_11111111_10010100_01011110_11101101_01101100_00010010_11111000_00110100_01101101_10101001_11111111_00001010_01111000_01000000_01111100_00000011_10101111_10001100_11010101;
assign in[270] = 496'b11111100_00001110_01100101_01001100_01011000_11111111_10000011_01000110_11100000_11111111_10010110_11111111_11111111_01011011_11000000_11111111_11111111_11111111_11111111_11111001_01111100_11110110_11111111_11111111_11111111_11111111_11111111_01011001_10100110_11001111_10101010_11001111_11111111_11111111_10111101_01001000_01110100_01100110_11000010_11111111_11111111_11111111_11100111_01110000_10111110_11111111_10111100_00000001_00001001_01101100_00100000_11111111_11111111_01100001_00110100_10000110_10010000_11111100_11111111_11111111_11111111_11111111;
assign in[271] = 496'b11111111_11101100_10100000_11110101_11111111_11111100_10011100_01000010_01110110_01010101_10111011_11101100_00001010_11011000_10000001_10010011_11100101_01001100_10100000_11110101_10001000_00100110_11111111_11100010_01001001_00100010_00100001_10000010_11111001_11111111_00010010_10000011_10101011_11010001_11111111_11111111_11000111_01010010_11101111_11111111_11111111_11111111_11011000_01011100_11000110_11111111_11111111_11111111_11101110_01010001_10011011_11111111_11111111_11111111_11111111_00100110_10010101_11111111_11111111_00011101_11111111_11111111;
assign in[272] = 496'b10001101_01110110_01111011_01111100_01110000_10001111_01111000_01010110_10010111_11101011_10011000_11000101_01100011_00101011_11110001_11111111_11111111_11110001_00011110_01101011_11011101_11111111_11111111_11111111_11110001_01100001_10100010_11111111_11111111_11111111_11111111_10110001_01111100_11000101_11111111_11111111_11111111_11111111_11011000_01001100_11111111_11111111_11111111_11111111_11001111_01110011_01001011_11011000_11100111_10010011_00101101_01110111_01001010_01110001_01111011_01111011_01111100_01100001_10000110_10000010_11000010_11111010;
assign in[273] = 496'b11111111_11111111_01000100_11001011_11111111_11111111_11111111_11111000_01100000_11101111_11111111_11111111_11111111_11111111_11000101_00110001_11111111_11111111_11111111_11111111_11111111_00010000_10011101_11111111_11111111_11111111_11111111_11100110_01001100_11101110_11100110_11101100_11111111_11111111_10110101_00010100_11111111_00101111_11010010_11111111_11111101_01001000_00011101_10110011_01001101_11111100_11111111_00000001_00111010_10111011_01001110_00000110_11111111_11100110_01100111_11011011_11111111_11010011_11101111_11111111_11111111_11111111;
assign in[274] = 496'b11111111_00001001_10011101_11111111_11111111_11111111_11111111_01001000_11011010_11111111_11111111_11111111_11111111_11101110_01010101_11111111_11111111_11111111_11111111_11111111_10111001_00110100_11111111_11111111_11111111_11111111_11111111_00011011_10110001_11110111_00111011_11111111_11111111_11110110_01011111_11111101_10001111_00111010_11111111_11111111_10100101_01100111_00101110_01101100_11010010_11111111_11111111_00100011_00100000_00011100_10100001_11111111_11111111_11111111_10101101_11111011_11011011_11111010_11111111_11111111_11111111_11111111;
assign in[275] = 496'b11111111_11111111_01000111_11100100_11111111_11111111_11111111_11100110_01001000_11111111_11111111_11111111_11111111_11111111_00001001_10011001_11111111_11111111_11111111_11111111_11110011_01100011_11111010_11111111_11111111_11111111_11111111_10010100_10001100_11111111_10110001_11000111_11111111_11111111_01010101_11101010_11111011_01011000_11010011_11111111_10100011_01111101_00000011_10001010_00100001_11111111_11110100_01010000_10111110_10001101_01101011_11100100_11111111_11100010_10111110_11111111_11111111_11000010_11111111_11111111_11111111_11111111;
assign in[276] = 496'b01101000_00011011_01100001_01011110_11111111_11111111_01111000_10001110_11100011_01010000_00010110_11111111_11111111_10001010_01111101_10011110_00110011_01001011_11111111_11101011_10000111_01110111_01111101_01101110_11010001_00100000_01101111_01111100_01110100_01001000_01110100_11110111_10010100_10000001_01111000_10101010_11100011_01101100_10000011_11111111_00010011_00101001_11111111_11111111_00010011_00111110_11111001_01100110_10101000_11111010_11000001_01010000_00001101_11101001_01111000_01011100_01100110_01011111_10001011_10001000_11000110_11111010;
assign in[277] = 496'b00010011_01110100_01111011_01101011_00011101_10011100_01100101_11000001_11110011_11011000_10100010_11111111_10010011_00001010_11111111_11111111_11111111_11111111_11111111_11111011_00101010_00010111_11010100_11111111_11111111_11111111_11111111_11111011_10010010_01011101_11111001_11111111_11111111_11111111_11111111_11011010_01011100_11001111_11111111_11111111_11111111_00001001_01111101_01000110_11111011_11111111_11111111_11000010_01111011_00011010_11111101_11101001_11111111_11111111_11010111_01110001_01101000_01000111_01100100_11101000_10010010_10000001;
assign in[278] = 496'b01011100_01111101_10111110_11111111_11111111_11110101_01100111_01111101_11000100_11111111_11111111_11111111_11110001_01101011_01111100_11010100_11111111_11111111_11111111_11111111_01011100_01111001_11110010_11111111_11111111_11111111_10110110_01111101_01001000_11111111_11111111_11111111_11111111_00100111_01111101_00110101_11111111_11110010_10111100_11111111_00111000_01111101_01110100_00101001_01011000_01111101_11111111_10000001_01111011_01111101_01111110_01111101_01111101_11111111_11111111_11011100_10110010_10100010_10110000_11111111_11111111_11111111;
assign in[279] = 496'b11111111_11111111_00100011_10010000_11111111_11111111_11111111_11101110_01110100_10101000_11111111_11111111_11111111_11111111_10011001_01111101_11110100_11111111_11111111_11111111_11111111_01001011_00111111_11111111_11111111_11111111_11111111_11111111_01111100_10000110_11111111_11111111_11111111_11111111_11011010_01111101_10101011_11111111_11111111_11111111_11111111_10010000_01111100_11100100_11111111_11111111_11111111_11111111_00001010_01011000_11111101_11111111_11111111_11111111_11111111_00101001_00101001_11111111_11111111_00011101_10001001_11111111;
assign in[280] = 496'b11111111_11111111_11111111_10001011_00100011_11111111_11111111_11111111_11100110_01100000_11001000_11111111_11111111_11111111_11111111_01000010_00001010_11111111_11111111_11111111_11111111_10110110_01011101_11111011_11111111_11111111_11111111_11111111_01010001_10101100_11111111_11111111_11111111_11111111_11001101_01101001_11111111_11111111_11111111_11111111_11111111_01000000_00010011_11111111_11111111_11111111_11111111_11010011_01100111_11101100_11111111_11111111_11111111_11111111_10100111_00100011_11111111_11111111_11111111_11000000_11111111_11111111;
assign in[281] = 496'b00011011_01110100_01111101_01011001_11110111_01110010_01110001_00001110_00100110_00100101_11111100_01100101_01011100_11100001_11111111_11111111_11111111_11111111_01111101_10110100_11111111_11111111_11111111_11111111_11111111_01100010_00000111_11100101_11111111_11111111_11110100_10110111_10111100_01001111_01111010_01011110_01011110_01101011_01111101_11111111_11111110_11010010_00111100_01111101_00101110_10010110_11111111_11111111_11111111_00011010_01011100_11111110_11111111_11111111_11111111_11111111_10010110_01101100_00001011_11111111_11111111_11000010;
assign in[282] = 496'b10101110_11111001_11111111_11111111_10101101_00000110_11111111_11111111_11111111_11111111_11111111_00110111_11010110_11111111_11111111_11111111_11111111_11111111_10101010_00100001_11111111_11111111_11111111_11111111_11111111_11111110_00110111_10011110_11111111_11111111_11111111_11010110_11111111_11110110_00101011_00010000_10110001_10011010_01011100_11111111_11111111_11111111_11000001_10000011_10001111_01101000_11111111_11111111_11110111_11110000_11000000_11000110_01011110_01001001_01001100_00111000_01001000_00111100_01001000_11111111_11111111_11111111;
assign in[283] = 496'b11111111_11111111_01010000_11101011_11111111_11111111_11111111_11101111_01101110_11111000_11111111_11111111_11111111_11111111_10111100_01100011_11111111_11111111_11111111_11111111_11111111_00010010_00001101_11111111_11111111_11111111_11111111_11111111_00110000_00000100_11111111_11111111_11111111_11111111_11111111_00111001_10011000_11111111_11111111_11111111_11111111_11110100_01111001_11010001_11111111_11111111_11111111_11111111_11110000_01110010_11111000_11111111_11111111_11111111_11111111_11101001_01101010_11111111_11111111_11110000_01100011_11111111;
assign in[284] = 496'b11010100_01000101_01001111_11100111_11111111_11111111_00100010_10101101_00011101_11001000_11111111_11111111_11111111_01010000_11100011_01011100_11111100_11111111_11111111_11111111_00011000_01001100_00010110_11111111_11111111_11111111_11111111_11001110_01111001_01001001_10100000_11111111_11111111_11111010_00110011_10101101_11010111_00101101_10110110_11111111_00001011_00001101_11111110_11111111_00000010_10110110_11000111_00111011_11111111_11111111_10110011_00111100_11111011_11001100_00111110_10111100_00011011_00100000_11110011_10001010_11001100_11111111;
assign in[285] = 496'b00000100_11111111_11111111_11111111_11111111_10111100_00000111_11111111_11111111_11111111_11111111_11111111_11111111_00010110_11111111_11111111_11111111_11111111_11111111_11111111_00101101_10011111_11010101_11101010_11000100_11111111_11111111_00011000_00001100_10011110_00000000_00111110_11111111_11111111_11011110_10001111_11111111_10011100_00011011_11111111_11111111_11001000_00011010_10101000_00011111_11110011_11111111_11111111_11111111_01011101_00000101_11011010_11111111_11111111_11111111_11000110_00110101_11111110_11111111_11111111_11111111_11111111;
assign in[286] = 496'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_10011100_01011011_11011000_11111111_11111111_11111000_00001001_10000101_01100000_00111100_11111111_11111111_10111101_11101111_00000011_10101101_00110101_11111111_11110101_11111110_10000111_10101001_10001110_10100001_11111111_10001001_10000110_11001010_11110101_01010100_11110010_11111111_11111111_11111111_11111111_10010010_10000010_11111111_11111111_11111111_11111111_11111110_00111111_11110111_11111111_11111111_11111111_11111111_11000011_00010111_11111111_11111111_10000100_10100101_11111111;
assign in[287] = 496'b11000000_10100001_11111111_11111111_11111111_11111111_10111001_10110101_11111111_11111111_11111111_11111111_11111111_11000100_10101001_11111111_11111111_11111111_11111111_11111111_10101101_11001001_11111111_11111111_11111111_11111111_11111111_10100001_11001100_10101001_10010101_11111111_11111111_11111111_00011111_00110011_10101100_00000000_11111100_11111111_11111111_10100001_10101001_11111111_10010101_11111111_11111111_11111111_10100001_11010100_11111111_00010000_11111111_11111111_11111111_10100001_11011000_11111111_10010000_11111111_11111111_11111111;
assign in[288] = 496'b11111111_00000001_10100100_11111111_11111111_11111111_11110100_01000111_11110001_11111111_11111111_11111111_11111111_10010011_10010101_11111111_11100101_11101000_11111111_11111001_01001100_11011000_00011100_00100011_01010001_11111111_10011101_01011110_00100000_11100011_11100010_01010011_11110010_01101010_10010011_11111111_11101011_01001010_10110011_00010101_00011001_11111111_11100011_01001101_10101000_11111111_00101010_01000000_10010111_01000100_11001011_11111111_11111111_11111111_10100111_10011100_11111001_11111111_11111111_11111111_11111111_11111111;
assign in[289] = 496'b11111111_11110001_00110011_11111111_11111111_11111111_11111111_11011000_01100101_11111111_11111111_11111111_11111111_11111111_10100110_01000101_11111111_11111111_11111111_11111111_11111111_00001101_00111001_11111111_11111111_11111111_11111111_11111111_00001101_10011111_11111111_11111111_11111111_11111111_11111111_01011001_11010001_11111111_11111111_11111111_11111111_11111111_01111101_11100100_11111111_11111111_11111111_11111111_11111111_01111110_11100100_11111111_11111111_11111111_11111111_11111111_01001100_11011110_11111111_11111111_00000001_10101011;
assign in[290] = 496'b11111111_10110010_01111010_11000011_11111111_11111111_10110110_01111011_00010011_11111111_11111111_11111111_11110111_01101000_00111000_11110100_11111111_11111111_11110101_00111010_01100001_11110100_11111111_11111111_11111111_00110111_01101001_10111011_11111111_11111111_11111111_11111111_01111100_10011100_11111111_11111111_11111111_11111111_11111111_01010100_11101100_11010100_10100010_00000110_00101101_01110111_01111011_01111100_01110000_01011101_00110110_00001110_10100011_10111101_10110011_11100010_11111111_11111111_11111111_11111111_11111111_11111111;
assign in[291] = 496'b11110110_01110000_00100111_01101100_00011100_11111111_10011011_00111001_11111111_11101010_10011100_11111111_11111111_00001011_00001011_11111111_11111111_11111111_11111111_11111111_10001101_00101010_11111111_11111111_11111111_11111111_11111111_11011011_01100111_11011010_11101010_11100010_11111111_11111111_11111111_10011101_01011110_01110111_00101101_11111111_11111111_11111111_11111111_10100000_01100110_11011111_10000001_10000010_10100011_11011010_01000100_11101011_11111111_00100011_00000101_00100111_10101001_10000101_11111111_11111111_11111111_11111111;
assign in[292] = 496'b01111000_00100110_10010100_10010100_11011001_10101001_01111010_00010000_11111110_11111111_11111111_11111111_11111111_00011000_01111110_00100011_11111111_11111111_11111111_11111111_11111011_10000100_01111010_01001001_11101110_11111111_11111111_11111111_11111111_10100110_01111101_00101101_11111111_11111111_11111111_11111111_11111111_10100001_01111100_11111111_11111111_11111111_11111111_11111111_11111001_01000100_00101111_00110100_00110100_01000100_01111100_00011111_01011101_00110101_00010001_10010100_10010011_10101101_00010001_11111111_11111111_11111111;
assign in[293] = 496'b00100100_01000010_01001000_00110101_10110001_00011101_11010110_11111111_11111111_10101000_11000010_00100011_11111111_11111111_11111111_11111111_11111111_11111111_01001101_11001000_11111111_11111111_11111111_11111111_11111111_11100010_01001010_00010100_11011010_11111111_11111111_11111111_11111111_11111001_10101100_00111000_01011001_01000110_00101001_11111111_11111111_11111111_11111111_00001111_00100000_11101110_11111111_11111111_11111111_11111101_01100011_11101100_00001001_11111111_11111111_11111111_11111100_01100011_10011010_11111111_11111111_00110010;
assign in[294] = 496'b11111111_11111111_00001101_10111011_11111111_11111111_11111111_11110101_01010010_11111111_11111111_11111111_11111111_11111111_10011000_10001010_11111111_11111111_11111111_11111111_11111010_01001101_11110001_11111111_11111111_11111111_11111111_10011111_00000000_11111111_11001100_00010101_11111111_11111010_01001101_10111001_11011011_01010011_10001110_11111111_10011110_01110100_00101000_01110011_01010011_11111010_11111111_01010001_10010110_11111111_10000011_11011011_11111111_11111111_10110011_11111111_11111111_11111111_11111111_11111111_11111111_11111111;
assign in[295] = 496'b11111111_11111111_11111111_11111111_11110000_11111111_11111111_11111111_11111111_10100000_01101111_11111111_11111111_11111111_11111111_00000000_01111111_01111111_11000000_11000000_10010001_01010000_01111111_00011111_11100000_01111111_01111111_01100000_01101111_01100000_11111111_11111111_11111111_11111111_11111111_00100000_00100000_11111111_11111111_11111111_11111111_11111111_01010000_10010001_11111111_11111111_11111111_11111111_11111111_01111111_11000000_11111111_11111111_11111111_11111111_11111111_01111111_11000000_11111111_11111111_00101111_01101111;
assign in[296] = 496'b11111110_01100111_11011011_11111111_11111111_11111111_11000101_01010111_11111111_11111111_11111111_11111111_11111111_10001100_10001011_11111111_11111111_11111111_11111111_11111111_00100001_11010111_11111111_11111111_11111111_11111111_11110101_01011111_11011000_11010101_10011000_11101000_11111111_10010110_01110111_01100101_00101100_00011111_00110011_11111010_01010100_00011011_00000011_11111111_11110110_01011111_11101111_00011100_11111001_00111100_10100111_00111000_00001100_11111111_11111111_11111111_10011101_10000110_10110111_11111111_11111111_11111111;
assign in[297] = 496'b11111111_11111111_11111111_11111111_11111111_11111110_10000100_01001001_01111101_01001100_11011111_11001111_01001010_01101001_01111101_00000111_01010110_00101010_01101010_00010011_10011111_01111101_11100001_10011100_01110101_00110111_10000111_01100111_10010001_11111110_10100000_01111001_01110111_00100110_10111000_11111111_11110110_01011100_00011001_11111111_11111111_11111111_11111111_10011001_01110001_11011001_11111111_11111111_11111111_11111000_01011101_10000011_11111111_11111111_11111111_11111111_00001001_01011110_11110110_10110000_01101101_11001101;
assign in[298] = 496'b00100000_00101011_11100000_11111111_11111111_11110111_01100111_01111101_10100110_11111111_11111111_11111111_11110100_01101100_01111101_10100110_11111100_10010101_10011111_11000110_01111101_01111101_00010100_00110011_01111101_01111011_01011000_01111101_01111101_01100000_01111011_01111101_00001001_01100001_01111101_00111000_11111101_01101000_01111101_11111010_01011110_01111101_00010011_11101111_01110001_01111101_10101010_01111101_01111101_10111100_11011000_01111101_01111101_00110010_00101111_10100110_11111111_11111111_01011110_11111111_11111111_11111111;
assign in[299] = 496'b01101000_01000000_00110000_01100100_00000010_00100000_10000110_11111111_11111111_11111011_00100011_11100110_01101001_11101110_11111111_11111111_11111111_11111001_11110111_01100110_11010100_11111111_11111111_11111111_11111111_11111111_10011001_01010010_11101011_11111111_11111111_11111110_11111111_11111111_10001001_01100000_10001000_00001000_01011101_11111111_11101101_11000110_11001001_10100110_10001110_01110110_00010110_01100010_01010100_01101000_00011001_00011001_00110010_00110010_11101110_11111111_11100110_01001010_01100011_11111111_11111111_11111101;
assign in[300] = 496'b11110000_11111111_11111111_11111111_11111111_01111111_11000000_11111111_11111111_11111111_11111111_11111111_01000000_10010001_11100000_11000000_11000000_11100000_11111111_00100000_01101111_01000000_01000000_01010000_01101111_11000000_01111111_10110000_11111111_11111111_11111111_10100000_01101111_01111111_11000000_11111111_11111111_11111111_11000000_01100000_01111111_11010000_11010000_11111111_10100000_01101111_11110000_10010001_01010000_01111111_01111111_01111111_01000000_11111111_11111111_00100000_11000000_11111111_11111111_11111111_11111111_11111111;
assign in[301] = 496'b01111000_00110110_10111010_11111111_11111111_01110100_10110001_11010011_00011111_00011100_11111111_10011101_01110110_11010110_11111111_11111001_01001111_11000000_11111110_10100000_01011010_00010100_11001010_00011001_00010101_11111111_11111111_11110011_10010011_00101001_00110111_00010010_11111111_11111111_11111111_11111111_10111001_01111110_10110101_11111111_11111111_11111111_11100110_01100010_01000101_11111111_11111111_11111111_11100110_01011001_01101100_11011100_11111111_11111111_11010011_01011000_01011100_11011001_11111111_01000000_11101110_11111111;
assign in[302] = 496'b10011101_00010111_01100111_00010111_10001001_00101010_10010000_10110011_10111001_10010011_00110010_01011011_10111000_11111111_11111111_11111111_11111111_11101100_01011010_10101111_11111111_11111111_11111111_11111111_11111111_11010001_10101010_10100111_11011000_11100000_10111010_11100101_11111111_11111111_10111111_01110011_01111101_01111100_11001100_11111111_11111111_11101011_01101111_00111110_10101111_11111111_11111111_11111111_10111000_00101011_11111111_11110111_10111100_11111111_11111111_10011101_00010111_11001010_10001100_11101111_00110110_01110101;
assign in[303] = 496'b01000101_01111101_01100111_00111100_00011001_01111101_01001111_00010000_00001001_00001101_01011001_01111101_10110001_11111111_11111111_11111111_11111111_10101010_01011101_11111011_11111111_11111111_11111111_11111111_11100010_01111000_11011001_11111111_11111111_11111111_11111110_11100001_01011010_00110000_10011100_00011100_01000011_01011111_01111100_11000101_01011101_01111101_01111101_01111100_01100110_00101010_11111111_10011000_01111101_10011001_11010110_11111111_11110110_11111111_11100010_01110111_00100110_00000011_00000001_10010111_01010101_01111110;
assign in[304] = 496'b11111111_11100011_10011011_00110100_01111100_11111111_11000101_01110111_01111100_01111101_01111100_11111111_11111111_11111111_11001010_01110110_01111101_00110101_11111111_11111111_11011100_01101001_01001111_00000001_01110111_11111111_10100100_01100111_01000001_11110010_11011111_01111101_00100000_01111100_01010101_11101100_11111111_10101111_01111100_01111101_00110010_11000110_11111111_11000000_01110000_00101011_10110110_11111100_11111110_10101100_01100100_01000000_11011101_00100110_11000001_00001101_01111100_00101010_11110010_01100001_10000110_11111010;
assign in[305] = 496'b11111111_11111111_11111111_00110111_10111111_11111111_11001001_00011100_01001110_01111110_10101010_11111111_10001110_01111101_00110101_01011101_01111111_11001101_11001110_01111001_01010100_01100000_01111110_01111110_11010001_10100000_01111110_01111110_01100101_01011001_01110111_11110001_11111010_11000110_10111011_11100001_01101100_01000011_11111111_11111111_11111111_11111110_10101110_01111110_10101100_11111111_11111111_11111111_11101011_01100110_01100010_11101011_11111111_11111111_11011011_00101100_01111110_10001111_11111111_01110100_00010111_11101100;
assign in[306] = 496'b11100011_10001100_10101001_11111111_11111111_11111110_11000000_00101001_01001110_11011010_11111111_11111111_11001111_01000011_01111110_01100011_01110110_11010100_11100001_01101100_01111100_10000101_10101110_01111101_11011011_11010010_00010010_10110100_11111111_10001000_01111110_11011101_11111111_11111111_11111111_11111111_00110111_01101100_11110010_11111111_11111111_11111111_11100000_01111110_00011111_11111111_11111111_11111111_11111001_00111011_01111100_11100000_11111111_11111111_11111111_00011010_01111110_10010001_11111111_01100101_00110010_11111111;
assign in[307] = 496'b11000110_01110110_01111011_11010111_11111111_11111111_00100110_01111101_00111101_11111111_11111111_11111111_11100100_01111011_01111101_10111000_11111111_11111111_11111111_00010111_01111100_01100110_11111111_11111111_11111111_11011100_01100111_01111101_10101010_11111111_11111111_11111111_00011010_01111101_01010000_11111110_11111111_11111111_11110000_01110001_01111101_10000100_11111111_11111111_11000100_01011110_01111100_01111101_01011001_01000110_01001100_01000101_01010011_11010000_10110111_10000010_10101010_11101011_11111111_11111111_11111111_11111111;
assign in[308] = 496'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11101110_11100011_10101011_01001000_00100101_00110100_01011101_01110011_01111101_01111101_01000000_00001001_01000101_01111101_01111101_00111101_10100101_11111111_11111111_10001011_01111101_00001101_11111111_11111111_11111111_11000011_01110101_00110101_11111101_11111111_11111111_11111111_01001010_01110000_11110100_11111111_11111111_11111111_11111111_00110001_01110100_11100101_11111111_11111111_11111111_11101100_00110101_01100000_01101100_00101001_00000101_11111110_10100010_00110001;
assign in[309] = 496'b11111111_11111111_11111111_11111111_11111111_11100110_11111111_11111111_11111111_11111111_11111111_01111010_01111101_01011100_01000011_00011110_00010011_00110100_11011101_11010001_10001000_10001001_00100110_01111110_01110110_11111111_11111111_11111111_11101011_01000100_01011111_11000110_11111111_11111111_11101100_01010001_01001011_11101100_11111111_11111111_11111111_10010101_01111011_11010110_11111111_11111111_11110001_11111110_01010000_01100101_11001001_11110111_11110001_11111110_11111111_11010000_00111000_01111110_01110110_11111111_11111111_11101110;
assign in[310] = 496'b11110110_10001000_01100110_01110000_01110111_11110110_01000100_01100100_11010000_00100110_01111101_11100011_01001000_01001001_11100111_11111111_00010000_01111101_01011011_00111001_11110100_11111111_11110010_00111000_01111101_01101111_11101101_11111111_11111111_11010101_01110110_01111101_00100111_11111111_11111111_11111111_11100001_01110110_01111101_00101110_11111111_11111111_11001101_00010100_01111101_01011110_01111100_11010010_11110001_01010010_01111101_01110011_10011101_01110100_01111000_01110001_01111011_00110001_11000100_10100110_11010000_11111111;
assign in[311] = 496'b11111111_11111111_10100010_01111100_00010011_11111111_11111111_11100111_01011011_01110111_11001011_11111111_11111111_11111111_00100101_01111101_10001001_11111111_11111111_11111111_11011011_01111101_01110001_11111010_11111111_11111111_11111111_00011100_01111100_00010011_11111111_11111111_11111111_11111010_01100001_01111101_10111000_11111111_11111111_11111111_10111001_01111101_01101010_11110000_11111111_11111111_11111111_10101100_01111110_01100100_11011110_11111111_11111111_11111111_00010010_01111101_00001010_11111111_11111111_01001011_11011011_11111111;
assign in[312] = 496'b11110001_00001010_01111001_01101111_00100111_11111111_00101001_01111100_00100001_00100100_01110001_11111111_10010111_01111101_10001001_11111110_11111111_11101000_11110111_01111000_00110101_11111111_11111111_11111111_11111111_11111111_01010000_00110010_11010110_10110001_10100110_11111111_11111111_11101010_01111100_01111100_01111101_01100111_11100110_11101001_01010110_01110111_00101111_11000000_11111010_11111111_00010101_01111101_11001110_11111111_11111111_11111111_11111111_10101110_01101010_01001001_00001100_10100111_11000001_10100011_00010100_00010100;
assign in[313] = 496'b10110110_11001001_11101100_11111101_11111111_01110111_01101101_01111101_01111110_01110000_00100111_01111110_10110101_11111111_11011101_10111111_00001101_01110100_00100110_00000001_11111111_11111111_11111111_11111111_11101110_11111111_11001101_10100101_11000000_11101010_11111111_11111111_11111111_11111111_10100100_01111110_01111100_10011111_11111111_11111111_10011011_01111011_01110001_10000111_11110101_11111111_11001100_01111110_00001101_11110101_11111111_11111111_11111111_11111011_01001010_01001100_00010111_10000011_00010110_11011011_11000101_10010111;
assign in[314] = 496'b11111111_11111111_10110011_01101000_11110000_11111111_11111111_11111001_01010000_01011100_11111100_11111111_11111111_11111111_10100001_01111101_10011100_11111111_11111111_11111111_11110011_01100001_01000001_11111111_11111111_11111111_11111111_10100100_01111110_11001110_11111111_11111111_11111111_11111111_00100011_01111110_11100110_11111111_11111111_11111111_11111111_01001111_01100111_11111111_11111111_11111111_11111111_11111110_01010110_00100000_11111111_11111000_11111111_11111111_11111010_01110001_00000000_11111111_11111111_01000110_00000011_11111111;
assign in[315] = 496'b01110011_01110011_11110100_11111111_11111111_11101001_01111100_01011110_11111111_11111111_11111111_11111111_10100110_01111110_00001111_11111111_11111111_11101110_11111111_00110001_01111101_11000100_11111111_11111111_01001100_11011011_01111001_01001100_11111111_11111111_11101101_01110010_00100001_01111110_10101100_11111111_11111111_10001010_01111110_01111001_01101110_11000111_11110100_11100110_01101111_01111110_00101101_00110101_01110111_01110011_01111110_01111110_01111110_11111111_11111111_11110101_11010010_11000001_01101110_11111111_11111111_11111111;
assign in[316] = 496'b11000001_01111110_00111111_11111111_11111111_11111111_10000110_01111110_10001110_11111111_11111111_11111111_11111111_01010000_01110101_11001100_11111000_11111111_11111111_11001000_01111100_01111010_01110011_01011111_11100000_11111111_00100100_01111101_01101111_00100010_01111110_10001000_11100000_01111101_01010010_11011111_11001011_01111110_10001100_11000100_00000101_11110100_11110101_01000010_01011011_11111010_10000111_01101100_10011100_01011010_01110110_11010000_11111111_11111011_00110000_01111011_01001011_11010000_11111111_11111111_11111111_11111111;
assign in[317] = 496'b00000011_01111101_01000110_11010110_11111111_01100001_01111100_01111101_01111100_01110101_10100111_01001101_01111101_01111101_00111110_10000010_01011001_01110100_01111101_01100100_01100010_01010111_10111010_00011000_01111100_01111110_00001101_11101110_00110111_01111101_01111110_01111101_01111101_00001101_11111111_11101000_01110100_01111101_01111100_01000000_01100100_11011000_00001110_01111100_01111101_01111010_11001101_01101101_01010111_01100001_01111101_01111110_00110000_11111111_11010111_00111111_01111101_01111100_01111101_11111110_10110010_10010000;
assign in[318] = 496'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_10111010_01000001_01110001_00001011_11111111_10101001_00001001_01111011_00110000_10111001_01110110_11111111_11100100_01001111_01001100_01100111_01011010_01111011_11111111_11101001_01111100_10110010_11111011_10111011_10111101_11111111_11100010_01111110_11011101_11111111_11111111_11111111_11111111_11100010_01111110_11101111_11111111_11111111_11111111_11111111_11101001_01111100_11011110_11111111_11111111_11111111_11111111_11111111_00111011_10101100_11111111_11111111_10001011_00101100_11111111;
assign in[319] = 496'b01111101_01101110_01111100_00100001_11111000_11110011_11110011_11110110_11110011_10011000_11011110_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11110100_11111111_11111111_11111111_11111111_11111111_11111111_10111000_11111111_11111111_11111111_11111111_11111111_11111111_10010101_11010101_11111111_11111111_11111111_01011010_11000111_11111111_00010000_10101000_11000111_00011110_01010101_00101101_11111111_11110100_10100011_00001110_00000100_11010101_00101101_11111111_11111111_11111111_11111111_11111111_11100011_01001000_00000101_00000101;
assign in[320] = 496'b11111111_11111111_11111111_11111111_11111111_00000011_01000111_01111101_01011110_00011101_11111101_01011110_01100000_01110010_00011001_10101100_01011110_00010000_01010111_01001111_01100000_00110011_11111111_11100011_01100001_11100000_00110010_01101111_00111100_11111111_11111010_01101110_11111111_11111111_11111111_11111111_11111111_10101010_01101010_11111111_11111111_11111111_11111111_11111111_01000100_00001100_11111111_11111111_11111111_11111111_10101001_01101001_11100101_11111111_11111111_11111010_00000000_01100100_10000111_11010001_01111101_01011000;
assign in[321] = 496'b11111111_11111111_11111111_00001000_00011110_11111111_11111111_11111111_11010101_01101110_11010011_11111111_11111111_11111111_11111111_00011011_01100011_11111111_11111111_11111111_11111111_11001100_01110000_10111010_11111111_11111111_11111111_11111111_00101101_01000111_11111111_11111111_11111111_11111111_10101101_01110010_10111101_11111111_11111111_11111111_11111111_00110010_00111100_11111111_11111111_11111111_11111111_11011110_01111010_10010011_11111111_11111111_11111111_11111111_00000101_01111101_10101111_11111111_11111111_10110000_11010101_11111001;
assign in[322] = 496'b11111101_01001111_10011011_11111111_11111111_11111111_10000111_00011000_11111111_11111111_11111111_11111111_10010011_01010010_11111010_11111111_11111111_11111111_11110100_01101100_11001010_11111111_11111111_11111111_11111111_10010010_00101001_11111111_11111111_11111111_11111111_11111111_10100111_01000010_11101101_11111111_11111111_11111111_11111111_11111001_00101011_01010000_11000010_11111101_11111111_11111111_11111111_11111111_11000001_01001001_01100000_00101001_00011100_11111111_11111111_11111111_11111111_11001110_10100001_11111111_11111111_11111111;
assign in[323] = 496'b11011110_01100101_01111000_10111011_11111111_11111111_00111101_11010001_01001000_10001111_11111111_11111111_10111001_00001101_11111111_01100001_10011001_11111111_11111111_00001100_11010001_00000101_01110110_11110001_11111111_11111111_00001100_01001000_01111100_01111101_10100110_11111111_11111111_10011001_01101011_01110010_00101000_00100110_11111111_11111111_00001100_10010110_11110111_11101010_11000110_11110010_11111111_10010000_10001100_11101111_11000000_01001101_10110000_11111111_11100110_01101001_01100000_01110100_10001111_11001110_10010100_11100010;
assign in[324] = 496'b11111111_11111111_11110000_01101100_11010000_11111111_11111111_11111111_00001111_01011100_11111010_11111111_11111111_11111111_11110010_01110101_00001110_11111111_11111111_11111111_11111111_10011110_01111110_11011111_11111111_11111111_11111111_11111111_01001011_01001000_11111111_11111111_11111111_11111111_11010110_01111110_10100110_11111111_11111111_11111111_11111111_10010111_01110111_11101111_11111111_11111111_11111111_11111111_00101100_01001110_11111111_11111111_11111111_11111111_11111111_01011010_10010011_11111111_11111111_01011110_11001110_11111111;
assign in[325] = 496'b11111111_11111111_11111111_11110000_01100001_11111111_11111111_11111111_11111111_00011110_01010000_11111111_11111111_11111111_11111111_10100100_01111001_10111101_11111111_11111111_11111111_11101100_01101110_10000010_11111111_11111111_11111111_11111110_00100000_01100110_11110110_11111111_11111111_11111111_11000111_01111000_10011001_11111111_11111111_11111111_11111011_01000010_00111000_11111001_11111111_11111111_11111111_10100111_01110111_11010011_11111111_11111111_11111111_11111011_01011111_10000111_11111111_11111111_11111111_11110010_11111111_11111111;
assign in[326] = 496'b11111111_11111111_10010010_10111001_11111111_11111111_11111111_10100110_01000101_01101101_10100111_11111111_11111111_11111100_01001010_10111100_00100000_10000111_11111111_11111111_00011011_00110100_11101100_01101000_10111001_11111111_10111011_00011101_11101101_00101100_00101010_11111110_11111111_11100001_11111111_10010101_01100011_11101111_11111111_11111111_11111111_11000100_01100111_10110111_11111111_11111111_11111111_11110100_01010110_10100101_11111111_11111111_11111111_11111111_00101001_00010000_11111111_11111110_10110100_11100101_11111111_11111110;
assign in[327] = 496'b10110101_01010011_10011001_01011001_11111111_11111111_00100000_10101001_11111010_01100110_11111111_11111111_11111111_10001100_10010011_11001000_01000000_11111111_11111111_11111111_11010101_01010101_01000011_10011100_11111111_11111111_11111111_11111111_00111001_01010111_11111111_11111111_11111111_11111111_10111001_01010110_01001011_11000011_11111111_11111111_10110111_01100110_11010010_10111101_00111100_11111111_00000011_01101101_11011100_11111111_11110111_01011100_11111111_10011111_01000011_10011110_10100011_00001111_00101100_10000001_10000001_10011101;
assign in[328] = 496'b01000010_01110100_01111101_01111101_01000101_00110000_10011100_11000000_11010110_10110100_01100101_10110011_11111111_11111111_11111111_11111111_11111111_11000111_11001100_11111111_11111111_11111111_11111111_11111111_11111111_01001000_11110100_11111111_11111111_11111111_11111111_11111111_01110111_00010100_11111111_11111111_11111111_11111111_11111111_10010110_01111100_11010101_11111111_11111111_11111111_11100000_11111111_01001000_01101000_10111111_11111111_11100000_01000011_11111111_11010011_01010101_01111000_00100100_01011110_11110110_10000110_01010000;
assign in[329] = 496'b10110011_10000001_10000100_11001110_11111111_00000000_01000001_10000101_00000011_01100111_10010111_10011110_00011000_11111110_11111111_11111111_11011001_01110111_01010110_11110000_11111111_11111111_11111111_11111111_01111110_00100111_11111111_11111111_11111111_11111111_11110111_01111110_00100100_11111111_11111111_11111111_11111111_10001101_00111010_00110011_11111111_11111111_11111111_11110101_01011011_10111010_01000011_00000111_11110101_11111111_00100000_00110110_11111111_11110000_00100010_01001000_10110101_01010110_11111011_11100110_01010100_11000110;
assign in[330] = 496'b11111111_11111111_11111010_11101110_11111111_11111111_11111010_00100001_01001100_00111010_00111011_11111111_11111111_10100101_00011101_11111111_11111111_11111101_11111111_11111111_10000010_10111111_11111111_11111111_11111111_11111111_11111111_11000101_00100100_10110001_10011110_11110111_11111111_11111111_11111111_11010111_01001111_00111011_11110011_11111111_11101110_11001001_00100000_00100000_11111100_11111111_01001010_00111010_00000111_10011001_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111;
assign in[331] = 496'b11111111_10010001_01111100_00011110_11111111_11111111_10010000_01111010_01111101_01111011_11101011_11111111_11111111_00110011_01111101_01111101_01101110_11110000_11111111_11111111_00110011_01111101_01111101_00001101_11111111_11111111_11111111_00110011_01111101_01111101_11001000_11111111_11111111_11111111_00110011_01111101_01011010_11111001_11111111_11111111_11101101_01101110_01111101_10010010_11111111_11111111_11111111_00001000_01111101_01111101_11000011_11111111_11111111_11111111_00111100_01111101_01011011_11100101_11111111_01011111_11001001_11111111;
assign in[332] = 496'b11111111_11111111_11111111_11001000_01000111_11111111_10011101_11001111_10001000_01100011_10011101_11111111_11111111_10101011_01111111_01101010_11001111_11111001_11111111_11111001_00111000_01101010_01100011_00100011_01011100_11111111_00110001_00111111_11111001_10111001_10001111_11100100_00000000_01010101_11111001_11111111_11111111_11111111_11111111_01110001_11001000_11111111_11111111_11111111_11111111_11111111_00111000_11111111_11001111_01011100_10111001_11111111_11111111_00000111_10011101_01101010_10001000_11111001_11111111_10100100_11111111_11111111;
assign in[333] = 496'b10100101_01111101_01000010_11111100_11111111_11001011_01110111_01101001_11100100_11111111_11111111_11111011_01000110_01111001_10110111_11111111_11111111_11111111_10110100_01111101_00110010_11111111_11111111_11111111_11111111_01001011_01111101_11000011_11111111_11111111_11111111_11111111_01111101_01010111_11101100_11010100_10010101_00011101_01011100_01111101_01111101_01111101_01111101_01111101_01101001_01000010_10001011_00010001_00010001_10001110_11001101_11110111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111;
assign in[334] = 496'b11111111_11111111_11111111_11111111_11111111_10011011_00110110_01100100_01101000_10111110_11111111_01110000_01111101_01101010_00111110_01111101_01011101_11111111_01110001_00011011_11111000_00010101_01111101_01111101_11001111_01001100_01010001_11001010_01100101_01111101_01111101_11001100_11011110_01010101_01111101_01011101_00010001_01111101_10100010_11111111_11110011_10100101_11101011_10000100_01111101_10110011_11111111_11111111_11111111_11111110_01001111_01111001_11011101_11111111_11111111_11111111_11010000_01111101_01011010_11111111_00101100_01111101;
assign in[335] = 496'b10000001_11000011_11111011_11111111_11101110_01100000_01010001_01111101_01001101_10001001_01110111_10001110_11111111_11111111_11010011_01111110_01111110_01111110_11111111_11111111_11111111_10000110_01100001_00111000_00001111_11111111_11111111_11000011_01111100_10111001_11111111_11111111_11111111_11111111_00111001_00111101_11111111_11111111_11111111_11111111_11110100_01110011_10011001_11101110_11110110_11111111_11111111_11100110_01111110_00100110_01111010_01010100_11111100_11111111_11101011_01111010_01111110_01111110_01010001_00101100_01111110_01111010;
assign in[336] = 496'b00010111_11111111_11111111_11111111_11111111_01011101_10000011_11111111_11111111_11111111_11111111_11111111_00011110_00011001_11111111_11100101_11101110_11111111_11111111_00100111_01101111_01011010_01111111_01100010_10111001_11111111_10110100_01111110_00000000_10101001_00000111_01101011_11111111_11001011_01111100_11011100_11111111_11000000_01110100_11111111_11001110_01111110_11010000_11111111_11111010_01111110_11111111_11111111_01111001_11010000_11111111_11111011_01001110_11111111_11111111_01101111_11111011_11111111_11111111_10100100_11111111_11111111;
assign in[337] = 496'b01010111_11110110_11111111_11111111_11111111_10011101_00010110_11111111_11111111_11111111_11111111_11111111_00100011_10011000_11111111_11111111_11111111_11111111_11111111_01011101_11110111_11111111_10110100_00100001_10101000_11111111_01101011_11010001_00110001_00111101_10100111_01100100_11111111_01000000_01100101_00101101_11111100_11100100_01100010_11111111_10111110_01111110_00111010_00001001_01100010_00111010_11111111_11111111_10100010_01110111_01111111_01000110_11010110_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111;
assign in[338] = 496'b00100110_10001000_11111111_11111111_11111111_11111111_00111111_10110010_11111111_11111111_11111111_11111111_11111111_01001111_11010000_11111111_11111111_11111111_11111111_11111111_01010101_10010001_00010001_10111111_11111111_11111111_11110111_01111000_10101001_11001011_01001010_11001000_11111111_11101110_01111010_11101001_11111111_11010101_00110101_11111111_10010101_01111011_11100100_11111111_11101110_01010100_11111111_10101111_01011111_11100101_11110000_00100101_00000011_11111111_11110101_00001101_01101010_01000101_00000101_11111111_11111111_11111111;
assign in[339] = 496'b10101111_01100100_11111011_11111111_11111111_11111111_11010111_01111110_11010111_11111111_11111111_11111111_11111111_11111111_01101101_10100010_11111111_11111111_11111111_11111111_11111111_01101101_10111111_11111111_11111111_11111111_11111111_11111111_01101110_11000001_11111111_11111111_11111111_11111111_11111111_01101101_10100010_11111111_11111111_11111111_11111111_11111111_01100001_10100010_11111111_11111111_11111111_11111111_11111111_01101101_10100010_11111111_11111111_11111111_11111111_11111111_01101101_10100111_11111111_11110000_01101110_11101010;
assign in[340] = 496'b10100001_11111111_11111111_11111111_11111111_11010101_10000100_11111111_11111111_11111111_11111111_11111111_11100100_00010011_11111111_11111111_11111111_11111110_11111111_11111111_01000001_11001000_00010110_00000000_00110110_11111111_11111111_01000100_11001100_11111110_11111111_10101000_11111111_11111111_00111111_11110000_11111111_11111111_00000001_11111111_11111111_00011110_11101011_11111111_11111111_00011101_11111111_11111111_00000011_11011100_11111111_11111111_11000101_11111111_11111111_00000001_10111001_11111111_11111111_11010001_11100111_11111111;
assign in[341] = 496'b11111111_10111000_01011001_01010111_01011100_11111111_11001101_01101101_10110111_11111111_11111011_11111111_11111111_00011000_10001010_11111111_11111111_11111111_11111111_11111111_00010101_10101101_11111111_11111111_11111111_11111111_11111111_11011110_01000101_00101101_00101100_00001010_11111111_11111111_11111111_11111111_11011111_01011111_10001110_11111111_11111111_11111111_11111110_00101111_00010001_11111111_11111111_11111111_11001000_00100111_01011000_11110011_11111111_00011100_01011011_00110101_01000011_11101100_11111111_11111111_11111111_11111111;
assign in[342] = 496'b11111111_11111111_00011000_11110011_11111111_11111111_11111111_11111110_00100111_11111011_11111111_11111111_11111111_11111111_11011010_00001010_11111111_11111111_11111111_11111111_11111111_00001101_10100001_11111111_11111111_11111111_11111111_11111111_01000111_11011001_11111111_11111111_11111111_11111111_10101011_01100001_11111111_11111111_11111111_11111111_11111111_10000010_10000111_11111111_11111111_11111111_11111111_11111111_00011101_10100110_11111111_11111111_11111111_11111111_11111111_00110111_11010100_11111111_11111111_11111111_11111111_11111111;
assign in[343] = 496'b11110011_00110100_01001111_00001001_01110000_11111101_00111110_00000101_11111101_11000001_01010000_11111101_00011011_10001001_11111111_11111111_00111101_10100000_10101000_00110100_11111111_10101010_00110100_01101101_11111110_00110110_11000011_10110010_01110110_01110101_01100101_11010110_01011001_10101010_01011011_00101011_00001010_01001101_11011100_10111001_01100001_10100001_00111001_11000110_01100110_11111111_11110101_01000110_10111010_00011010_00111101_10001010_11111111_11100110_01010011_01001000_10001011_01000101_11111100_10000001_10000001_11011111;
assign in[344] = 496'b10111111_11111111_11101111_10000101_11010000_10000010_00111101_11110010_01001101_00010000_00011110_11111111_10000010_01001001_00101000_01000010_00011100_01001001_11111111_10110001_01111100_01111101_01100011_00001100_11111001_11111111_11110010_01101010_00111000_11001001_11111111_11111111_11111111_10000010_00111011_11111110_11111111_11111111_11111111_11101011_01110011_11010101_11111111_11001001_01010000_10111111_11001101_00101011_11111001_10001111_01110101_01011001_11100110_10111100_01100000_01001101_01111110_01100101_11001101_01000011_00101000_11011101;
assign in[345] = 496'b11111111_11111111_11111111_11111111_11111111_11011000_01001100_01111011_01101100_01011001_00111101_00001101_11000001_10100100_01000010_11111111_11111111_00010001_11011100_11101100_01010011_10101110_11111111_11111111_10011110_00111001_01111100_10001011_11111111_11111111_11111111_00010101_01111101_00000010_11111101_11111111_11111111_11110010_01110101_11101001_11111111_11111111_11111111_11111111_00010111_00101001_11111111_11111111_11111111_11111111_11001111_01100101_11101110_11111111_11111111_11111111_11111011_00111100_10110011_11111111_00000110_00011001;
assign in[346] = 496'b11111111_11111111_10101001_00101000_11111111_11111111_11111111_11110110_01011000_11100110_11111111_11111111_11111111_11111111_00010111_10000110_11111111_11111111_11111111_11111111_11000000_01011001_11110110_11111111_11111111_11111111_11111111_01010101_10110110_11111111_11111011_11111111_11111111_10000100_10000110_11111111_11010111_01100010_11100011_11101100_01011001_11111001_11101001_00111010_01101111_11110001_10101100_01011110_10001001_01001000_00101010_10110110_11111111_11111111_11101110_10001101_11000100_11111111_11111111_11111111_11111111_11111111;
assign in[347] = 496'b11110100_01011101_11010111_10100111_11110011_11111111_10110100_01000110_11111111_11111111_11111111_11111111_11111111_10110100_00011101_11111111_11111111_11111111_11111111_11111111_10010000_00110011_11110100_11111111_11111111_11111111_11111111_00001010_01111101_01100010_11001110_11111111_11111111_11111111_01101101_01010010_00010110_01010001_11111111_11111111_11111111_01110001_10101000_10101001_01100110_11111111_11111111_11111111_01011100_00010110_00001010_00111101_11111111_11111111_11111111_11100101_01010111_01101010_10101001_11111111_11111111_11111111;
assign in[348] = 496'b00111011_11111111_11111111_11010111_00101101_11101100_01110011_11101110_10010000_01110111_01111101_11111111_11111111_01000010_01011001_01111000_01111000_00100001_11111111_11111111_10100101_01110101_00111110_11001110_11111111_11111111_11010000_01011111_11001000_11111111_11111111_11111111_11110001_01010000_10011101_11111111_11101110_10001000_01010000_00010011_00000111_11111111_10101110_01011111_01111100_01000101_01000111_11101111_00011011_00111010_10000001_01110010_11011001_10001111_00110011_10011010_00100000_01010000_11001011_11010100_10010100_11110101;
assign in[349] = 496'b11111111_11111111_11100000_00101001_11111111_11111111_11111111_11111111_01000001_11000111_11111111_11111111_11111111_11111111_11001000_01001000_11001100_10011010_11111111_11111111_11011100_01000101_01001111_00111111_01000111_11010000_00011000_00110100_01000100_11111110_11101000_01010111_11111111_11111001_01000111_11011101_11111011_01000101_10101111_11111111_10111010_00100010_11111111_10110110_00001100_11111111_11111111_01000110_11001001_11111111_11111110_11101111_11111111_10100000_00100000_11111111_11111111_11111111_11111111_11111111_11111111_11111111;
assign in[350] = 496'b11111111_11111111_11111111_11111111_11111111_11001110_00110110_01010100_01010110_00101000_11001011_10110010_01110111_00100100_01101001_10101000_10001100_01100110_01110101_10110001_11110000_01011001_11110101_11111111_00110010_01101111_00111111_01000101_00010001_11111111_11111111_00110110_10100011_01001110_10010111_11111101_11111111_11110110_01100110_11111111_11111111_11111111_11111111_11111111_10011010_00110101_11111111_11111111_11111111_11111111_11110100_01011100_11010110_11111111_11111111_11111111_11111111_00010000_00110010_11111111_11000110_01101110;
assign in[351] = 496'b11111111_11111111_11100100_01010011_11100110_11111111_11111111_11111001_01000100_11000011_11111111_11111111_11111111_11111111_00101010_10011111_11111111_11111111_11111111_11111111_00000001_00001001_11111111_11111111_11111111_11111111_10011000_00011010_11111111_11111111_11111111_11111111_11000100_00101100_11111101_11111111_11100010_00100011_11011100_01000011_11101100_11111111_10101110_01101110_01110100_11100001_01001000_00111000_00110111_00101100_01010101_10011000_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111;
assign in[352] = 496'b11101011_01101101_01111101_01111101_01100010_11111111_11011110_01110111_10100101_11101100_11101110_11111111_11111111_11111111_00100000_01000000_11111100_11111111_11111111_11111111_11111111_11010110_01111100_10111010_11111111_11111111_11111111_11111111_11100001_01011101_00000100_11111111_11111111_11111111_11000001_01011011_00111100_11100101_11111111_11111111_10100010_01111001_00010111_11111011_11111111_11111111_11111111_01011010_00110110_11111111_11110001_11111111_11111111_11111111_01011111_01101111_01001111_01110100_00101000_11000100_10110010_11000100;
assign in[353] = 496'b11111111_11111111_11111111_11111111_11111111_01111100_01111100_01010110_10100110_11110100_11111111_01111100_01110111_01100101_01111100_01111100_00110000_11111111_01101011_01111001_00100110_01100100_01111100_01110101_11001001_11001100_01100101_01111000_01100111_01101000_01111100_00110010_11111111_11111001_10111010_11111111_11110110_01111100_01111100_11111111_11111111_11111111_11111111_11010000_01111100_01000001_11111111_11111111_11111111_11111111_10000011_01111011_10000111_11111111_11111111_11111111_11001011_01110100_00111111_11111111_00101000_01010100;
assign in[354] = 496'b01101001_11110001_11111111_11111111_11111111_00000111_01111010_11011001_11111111_11111111_11111111_11111111_11010100_01101110_01100000_11011000_11111111_11111111_11111111_11111111_10111100_01011001_01111110_00110111_11010010_11111111_11111111_11111111_11111100_10100001_01111001_01000100_11111111_11111111_11111111_11111111_11101111_01111000_10010000_11001011_10100001_10011001_00000001_00101110_01110111_11101100_00100111_01110110_01111000_01111110_01111110_00001000_11111111_11111111_11110111_11110111_00110101_01011101_11111001_11111111_10111001_11100000;
assign in[355] = 496'b10111101_01110100_01111100_01111100_00001001_11010110_01100100_01111110_01111101_01111101_01111001_11111111_10000010_01111100_01011010_11010100_10010011_01111100_11111111_10000010_01111101_01110010_10011010_11001010_01111101_11111111_11101000_01100111_01111101_01111011_00100000_01001101_11111111_11111111_11101000_01000100_01111101_01111101_10110101_00100010_00100010_00100010_00001100_01111100_01111100_00000100_01111100_01111101_01111100_01111101_01111100_01111100_10110101_11101110_11000000_01111011_01111101_01110110_10000001_10001011_10100101_11011101;
assign in[356] = 496'b11111111_11111111_00001000_10101111_11111111_11111111_11111111_11011111_00111110_11111100_11111111_11111111_11111111_11111111_00110011_11010001_11111111_11111111_11111111_11111111_11000100_00110010_11001101_11100101_11111111_11111111_11111111_01011010_01010001_01001101_01000001_11111111_11111111_10110101_01000000_11011111_11110001_00110000_11111111_11111111_00110011_11100001_11111100_00101011_10111111_11111111_11111100_01011100_11001000_01010111_10110000_11111111_11111111_11111111_00110110_01100010_10110111_11111111_11111111_11111111_11111111_11111111;
assign in[357] = 496'b11111111_11100010_10101011_10000111_10010000_00011110_01001101_01111110_01000100_10110001_10011101_10100001_01101101_10010111_10111100_00111000_00100101_11110111_01000111_11010001_11111111_11111111_11111011_10000110_01000011_00100000_11111111_11111111_11111111_11111111_11111111_11101111_10001101_11111111_11111111_11111111_11111111_11111111_11111111_10001100_11111111_11111111_11111111_11111111_11111111_11111111_01010001_11110100_11111111_11111111_11111111_11111111_11111111_00010001_01000001_11110111_11111111_11111110_00101100_00111100_11000101_10101010;
assign in[358] = 496'b01111101_01110110_00100110_11011101_11111111_10111111_11110000_10111001_01011111_10001001_11111111_01001101_11111111_11111111_11111111_11100101_11111111_11111111_01110110_11010111_11111111_11111111_11111101_10100111_11111001_00001000_01010000_10011001_11011000_00011000_01111101_10011101_11111010_10101000_01011110_01100100_00100110_00100100_00110011_11111111_11111111_11111111_11111111_11111111_11010110_01101011_11111111_11111111_11111111_11111111_11111111_11101101_01111101_11111111_11111111_11000111_00110001_01001001_01011010_01111110_00101100_10010101;
assign in[359] = 496'b11111111_11111111_11000011_01000110_11111000_11111111_11111111_11110001_01010100_10110111_11111111_11111111_11111111_11111111_00011000_00001011_11111111_11111111_11111111_11111111_11001010_01011000_11111100_11111111_11111111_11111111_11110110_00110011_11010000_11111100_10001000_11110000_11111111_10001000_10001001_11111111_10011101_01001110_11111111_11011110_01001111_11111010_10110100_01101101_11010100_11111111_00100000_01001110_00000010_01010110_10111111_11111111_11111111_10011111_10100010_10000011_11011000_11111111_11111111_11111111_11111111_11111111;
assign in[360] = 496'b11111111_11111111_10110011_01101100_01111100_11111111_11111111_10100000_01011111_10110000_00001010_11111111_11111101_10010100_01111001_11100010_11111110_00011111_11111111_00111101_01111100_01111101_01001011_01001101_01000111_11111111_00101001_00100011_11101111_11101111_11100011_11111010_11111110_01011001_10111110_11111111_11111111_11111111_11111111_11111010_01101001_10111110_11111111_11100101_11111110_11111111_11111000_01110010_10110001_10111000_01111100_10111001_11111111_11111111_00001000_01010010_00101100_01101000_11011100_10011110_10000001_11011101;
assign in[361] = 496'b11111111_11111111_11111111_00000000_10100011_11111111_11111111_11111111_11110011_01010101_11111100_11111111_11111111_11111111_11111111_10001011_00010011_11111111_11111111_11111111_11111111_11101100_01011000_11100101_11111111_11111111_11111111_11111111_10000011_00000100_11111111_11111111_11111111_11111111_11001001_01101101_11001101_11111111_11111111_11111111_11111111_00110100_10101100_11111111_11111111_11111111_11111111_10011010_00100101_11111111_11111111_11111111_11111111_10011101_00111011_11111001_11111111_11111111_11111111_11111111_11111111_11111111;
assign in[362] = 496'b11001010_11111111_11111111_11111101_11111111_11101011_11111111_11111111_11111111_11111111_11111111_00100010_10111010_11111111_11111111_11111111_11111111_11111111_11000110_00110111_11000000_11110001_11111110_11111111_11111111_11111111_11110111_10100101_00100111_00011110_01001000_01100001_11111111_11111111_11111111_11100010_00000101_01101001_01001001_11011001_10010100_01001100_01100001_10101000_11011011_11111111_01111101_01001111_00111100_01111001_01100100_01111101_10011100_01001001_01110001_01110100_01100100_01000110_00010011_11111111_11111111_11111111;
assign in[363] = 496'b01110011_01111101_01111100_01111101_10001111_01111101_01111101_00100100_11010010_00100000_01011110_01110001_01101010_11011101_11111111_11111111_11101101_01010011_01111011_01010101_11111011_11111111_11000001_00011010_10100011_00100000_01111101_01011011_00110001_01101010_01111110_01010011_11111100_00010111_01111100_01111101_01110010_00111010_11100001_11111111_10001000_01111101_00010100_11100110_11111111_11111111_11100001_01111100_00110110_11010110_11001111_00000100_01101001_11100101_01110101_01111100_01111101_01111100_01111001_10001001_10000001_10110000;
assign in[364] = 496'b11111111_11010001_10000001_10000111_11101011_11101011_00000011_10110111_00110111_11010110_00011011_11101111_00001010_11110010_11011010_00011110_11110101_00100111_10010000_10001110_10000101_00101011_11101101_10101111_10000011_11101000_00101111_00101000_11110001_11111111_00111101_11110000_11111111_11111111_11111111_11111111_10000010_10000100_11111111_11111111_11111111_11111011_10110110_01000111_11111110_11111111_11111111_11111111_11010111_01001101_11010001_11111111_11111111_11111111_11011011_01000000_11011011_11111111_11111111_11100110_11111111_11111111;
assign in[365] = 496'b00101111_00110000_00101111_10111111_11111111_11000100_01111011_01111100_01111011_01110010_11111111_11111111_10111001_01111010_01111011_01111010_01011101_11111111_11111111_11111111_01111011_01111100_01111011_00100001_11111111_11111111_11000100_01111010_01111011_01111010_01111011_00011011_00010001_01110111_01111011_01000000_00010111_01111100_01111011_01111010_01011101_10001000_00000011_00111110_01111011_01111010_10010110_11001000_01110001_01111100_01110111_01100100_10010110_11111111_11111111_00110000_10100000_11000100_11111111_11111111_11111111_11111111;
assign in[366] = 496'b01010101_01101001_00001001_00111100_01100110_01000001_01010110_11010001_11111111_11111111_11100000_11001000_01111101_10011111_11111111_11111111_11111111_11111111_00101010_01110101_11101010_11111111_11111111_11111111_11111111_00101000_01111001_10010100_10101110_10101110_10101110_10101110_11010001_01010001_01111101_01111101_01111101_01111101_01111101_11111111_11111011_11110011_11110011_11110011_00011110_01111101_11111111_11010111_11001000_11001000_10010000_01110000_00011000_01001011_01110101_01111101_01111101_01111101_01001011_10000001_10000001_10000001;
assign in[367] = 496'b11111111_11111001_10010000_01100111_01110110_11111111_11001011_01001010_00000100_11010000_11101001_11111111_10100100_00111001_11011101_11111111_11111111_00000111_11001001_01001010_11110001_11111111_11111111_11001010_01011111_00111100_11010110_11111111_11111111_11110100_01010100_10100111_00010000_11111111_11111111_11110001_00111000_10001010_11111111_10010100_11111111_11111111_00000110_00011101_11111111_11111111_10010100_11111111_11001011_01011100_11110111_11111111_11111111_00011111_10110000_01011011_10111010_11111111_11111111_11000010_11111111_11111111;
assign in[368] = 496'b11111111_01011101_11001111_11111111_11111111_11111111_11111111_01010010_11101000_11111111_11111111_11111111_11111111_11111111_01101100_11111111_11111111_11111111_11111111_11111111_11011011_00100111_11110101_11010011_11111111_11111111_11111111_10011110_10000110_00110000_00100100_00000001_11111111_11111111_00011001_00110110_11111001_11101001_00100011_11111111_11011101_01010000_11110110_11111111_00000010_10101100_11111111_10101011_10111000_11111111_10011000_00010001_11111111_11111111_11100001_01000010_00100111_00010101_11111111_11111111_11111111_11111111;
assign in[369] = 496'b11111111_11111111_11111111_00111000_11101011_11111111_11111111_11111111_10110010_00001110_11111111_11111111_11111111_11111111_11111111_01000111_11011101_11111111_11111111_11111111_11111111_11010110_00111000_11111111_11111111_11111111_11111111_11111111_00011100_10110010_11111111_11111111_11111111_11111111_11111001_01011100_11110010_11111111_11111111_11111111_11111111_10011101_00011100_11111111_11111111_11111111_11111111_11111111_00111000_11001000_11111111_11111111_11111111_11111111_11101011_01000000_11111111_11111111_11111111_10110010_11111111_11111111;
assign in[370] = 496'b00100000_10100011_11010111_00011001_10001111_01011010_11010011_11111111_11111111_11101100_01100001_00001111_10010011_11111111_11111111_11111111_11101100_01101010_00001111_10011010_11111111_11111111_11111111_11101100_01110011_00101010_10011010_11111111_11111111_11111111_11101100_01111101_01000010_00001000_11111111_11111111_11111111_00000101_01101010_11000101_01110101_11101101_11111111_11111000_01101010_01000000_11111111_01100000_10100010_11111111_10001010_01111011_10110101_11111111_00001011_01000011_00101101_01110000_10000111_10000101_11010010_11100100;
assign in[371] = 496'b11111111_11010111_01000010_01111101_01011101_11111000_00001110_01111100_01100000_00010100_00101110_11111111_00110001_01111101_00110000_11111001_11111111_11111111_11111111_01000110_01000100_11111100_11111111_11111111_11111111_11111011_01101010_11011011_11111111_11111111_11111111_11111111_11111111_00110010_01000000_11100001_11100011_11101100_11111111_11111111_11100010_01101010_01111101_01111110_01101111_10100001_11111111_10101101_01111011_00101101_01100000_00100100_10111010_11111111_00011100_01001011_11111110_11111111_11111111_01110110_11111001_11111111;
assign in[372] = 496'b11111111_11010001_11000101_11000011_00011011_11111111_11001110_00011011_11111111_11111111_11110010_11111111_11111111_00100101_11101001_11111111_11111111_11111111_11111111_11111111_00101110_11111111_10110001_00110000_00000010_11111111_11111111_10001101_10011011_11010001_00011000_11001111_11111111_11111111_11111111_11111111_10010110_10011000_11111111_11111111_11111100_10100100_00101100_00011001_11111111_11111111_00100110_00111010_01001011_10110101_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111;
assign in[373] = 496'b11111111_11110010_10010110_01110001_01000001_11111111_11111111_00001100_01011110_01000110_01111101_11111111_11111111_10010110_01110000_11011110_00101001_01101011_11000011_11111000_01010111_00000110_11111111_00101101_00011000_01010001_01001110_01111101_00001111_00110001_01101000_11011110_11100111_01100001_01101101_00011011_10001011_11110011_11111111_11111111_01110101_00100110_11111111_11111111_11111111_11111111_11101001_01111010_00101011_11111111_11111111_11001101_11101010_11111111_01010011_01101100_11000011_10011101_01110110_00111111_01111110_01000100;
assign in[374] = 496'b00100100_11111111_11111111_11111111_11111111_00100100_01111101_00100001_11001000_11111110_11111111_11111111_11111100_10100110_01011000_01111110_00111111_11100111_11111111_11111111_11111111_11111111_10111101_01111000_00011011_11111111_11111111_11111111_11111111_11101011_01111100_10010111_11111111_11111111_11111111_11111111_10110011_01111110_11010010_10110000_10111001_10100100_00010111_01101101_01111110_11101011_01100110_01100111_01001001_00000110_01100000_01001011_11111111_11111111_11111111_11111111_11111111_01110001_10011001_11111111_11111111_11111111;
assign in[375] = 496'b11111111_11110101_10111110_10010010_11111010_11111111_11000110_01001001_00101001_00110011_00011000_11111111_10111100_00100100_11101100_11111111_00110100_00110110_11100110_00110101_11111101_11110111_10000101_01111110_10001010_10000101_00100110_00101001_01110010_01100001_01100010_11101101_11101011_00101001_01011010_00011011_01011001_10111101_11111111_11111111_11111111_11111111_00010100_00001110_11111111_11111111_11111111_11111111_11000111_01000100_11111001_11111111_11111111_11111111_11101111_01010100_10111110_11111111_11111111_10110100_11111111_11111111;
assign in[376] = 496'b01010001_01101111_00110101_01100010_10010001_01011011_10100110_11111010_11111111_11001101_01110011_01101100_11010101_11111111_11111111_11111111_11111111_00011101_00010110_11111111_11111111_11111111_11111111_11111111_10011011_00011000_11111111_11111111_11111111_11111111_11111111_00100111_01100111_11110101_11111111_11111111_11111111_11111111_01001001_01101010_00001101_11111111_11111111_11111111_11100100_01110010_10100100_01111010_00011101_11000000_11111110_00100010_00011101_11111111_10010111_01101000_01111110_01001101_01011010_11101010_10010111_10010101;
assign in[377] = 496'b11110110_11000111_10110011_10110011_10110011_01101010_01110000_01111110_01011111_01111101_01111110_11011000_10101001_11010110_11101101_00110100_01011010_11000000_11111111_11111111_11111111_00001011_01101010_11101000_11111111_11111111_11111111_11011010_01101111_10111010_11111111_11111111_11111111_11111111_00111101_00100110_11111111_11111111_11111111_11111111_11010101_01111100_11011100_11111111_11111111_11111111_11111111_10110011_01011000_11111111_11111111_11111111_11111111_11111111_11010111_01111001_11100000_11111111_11111111_00011001_01011110_00100111;
assign in[378] = 496'b10111010_11010001_10010101_10000010_10101100_00100010_01111010_01111110_01101101_00101110_10100101_11111111_11111111_11110111_01110101_10111000_11111111_11111111_11111111_11111111_11110000_01111000_11011011_11111111_11111111_11111111_11111111_11011001_01111110_11111111_11111111_11111111_11111111_11111111_11010100_01100110_11111111_11111111_11111111_11111111_11111111_00000010_01001011_10011100_01010101_10101101_11111111_11111111_00111001_01111110_01001001_00101101_11011101_11111111_11100011_01110110_00100010_11111111_11111111_01100000_11110101_11111111;
assign in[379] = 496'b11111111_11111111_11011010_01111100_01010000_11111111_11111111_11111111_01001100_01111100_10101011_11111111_11111111_11111111_10110110_01111100_00101011_11111111_11111111_11111111_11111111_01001101_01110111_11001010_11111111_11111111_11111111_10101101_01111010_01001010_11111111_11111111_11111111_11111111_00101011_01111101_10111110_11111111_11111111_11111111_11111111_01000000_01111101_11111111_11111111_11111111_11111111_11011101_01100111_10010011_11111111_11111111_11111111_11111111_00010001_01111100_11100010_11111111_11111111_01011010_11101011_11111111;
assign in[380] = 496'b11111101_01110001_11110001_11111111_11111111_11111111_11011010_01110101_11111111_11111111_11111111_11111111_11111111_10100100_00110011_11111111_11111111_11111111_11111111_11111111_00010101_10001000_11111111_11111111_11111111_11111111_11111111_01010010_11100101_11111111_11111111_00111001_11111111_11100110_01100001_11111010_11111111_11111111_01000111_11111111_10100001_00011101_11111111_11111111_11100110_01001101_11111111_00110100_01000100_10010001_10010010_00011001_00011011_11111111_10110011_10011001_10000001_10000001_10011001_11111111_11111111_11111111;
assign in[381] = 496'b11111111_11011001_10111101_10011011_10111100_11000000_01001001_01011101_00110100_00110100_01110100_10110011_01100100_10110110_11111110_11111111_11111111_01100111_01011011_11001101_11111111_11111111_11111111_11011001_01101101_01100111_11111111_11111111_11111111_11111111_01001010_00000110_01011000_11111111_11111111_11111111_11011110_01110010_11110001_00101011_10111010_11111111_11111111_00010100_00101001_11111111_11100000_01010010_11111110_11011101_01101000_11100000_11111111_11111111_00101100_10001101_00001111_00001001_11111111_01101011_01111001_11110001;
assign in[382] = 496'b01001110_01000100_01110001_11010000_11111111_00111010_11111110_11111110_00101010_00011001_11111111_01011010_11010101_11111111_11111111_10111110_01010101_11111111_01001100_11111111_11111111_11111111_11100111_01110110_11101110_00111010_11111111_11111111_11111111_11100111_01111101_11100111_01010011_11110100_11111111_11111111_11111110_01100111_11100111_00100010_00000100_11111111_11111111_11111001_01101100_10000100_11100100_01011010_10011011_11111110_11100010_01110011_01001011_11111111_11010000_01001110_01000011_00111110_01111011_11111001_10101010_10000001;
assign in[383] = 496'b11111111_11110011_10100101_10001000_11001101_11111111_10111110_01101000_00111100_00100100_01110010_11111111_11010010_01100111_10111100_11111111_11111111_00100110_11111111_00111010_10010111_11111111_11111111_11100100_01110110_11010010_01001001_11111111_11111111_11111111_00011011_00101110_11000010_00100001_11111111_11111111_11001001_01110011_11011000_10101011_00110001_11111111_11111100_01000010_10000010_11111111_11110000_01010111_11111011_10000101_00100111_11111111_11111111_11111111_01000101_00010100_01011010_11100010_11111111_01111101_10001111_11111111;
assign in[384] = 496'b10101000_01000000_01111011_01110010_00011010_00011101_01010111_10101101_11011010_11000011_01111001_00000001_01001010_11110011_11111111_11111111_11111111_01110100_01100100_11100011_11111111_11111111_11111111_11100000_01111100_01001010_11111111_11111111_11111111_11111111_10110100_01110000_01111010_10101111_11111111_11111111_11111111_00100000_01101001_01101111_10111011_11111111_11111111_11111111_01001111_10000110_10101000_01011010_11101110_11111111_10011010_01011110_11110010_11111111_00011101_01011110_10001010_01100100_11010000_10110101_01011111_10010000;
assign in[385] = 496'b11111111_11111111_01010101_10101011_11111111_11111111_11111111_11101011_01111000_11101011_11111111_11111111_11111111_11111111_10001111_00110001_11111111_11111111_11111111_11111111_11111111_01010101_10101011_11111111_11111111_11111111_11111111_10110010_01111111_11111001_11111111_11111111_11111111_11111111_00010101_01011100_11110010_11111111_11111111_11111111_11111111_00111000_10010110_11111111_11111111_11111111_11111111_11110010_01111111_11001000_11111111_11111111_11111111_11111111_11110010_01111111_11101011_11111111_11111111_10001111_11111111_11111111;
assign in[386] = 496'b00010111_01001110_00101101_00000010_00000010_00110111_00011101_11110010_11111111_11111111_11111111_11101111_01111101_11100110_11111111_11111111_11111111_11111111_11110101_01110110_10111110_11111111_11111111_11111111_11111111_11111111_00100110_01001101_10010110_00010011_10011110_11111111_11111111_11011110_01111011_01001101_10000110_11010000_11111111_11111111_10000100_01001101_11111111_11111111_11111111_11101101_11111111_01000101_10101000_11111111_11111111_11101101_00011110_11111111_00101011_00101011_10001110_00000001_01011000_10010111_10000001_10011000;
assign in[387] = 496'b10000001_10001001_11011111_11111101_11111111_01111101_01101000_01010011_01111101_00000101_11111110_01111101_01101100_11100010_11111000_01101101_01111101_10101101_01111101_01000011_10111000_00000111_01110110_01111101_00101011_00001011_01001001_01111001_01101101_01111101_01111101_00110001_11111111_11111111_11110010_11101101_01110000_01111110_10000010_11111111_11111111_11111111_10000011_01111101_01111101_11000000_11111111_11111111_11111111_01010010_01111101_00111011_11111111_11111111_11111111_11001101_01101011_01111101_10101010_01100101_01111101_01011011;
assign in[388] = 496'b11111111_11111111_11101111_00000000_10101100_01110000_00111001_11011111_00111110_01111001_01100001_11001000_10101100_00110110_01111101_01111101_01011010_00011011_11111111_11111111_11111100_01000010_00111001_10001000_11111000_11111111_11111111_11000110_01111101_11100100_11111111_11111111_11111111_11111111_00011000_00110011_11111111_11111111_11111111_11111111_11110111_01100000_10011111_11111111_11111111_11111001_11111111_11101100_01110010_10111010_11111111_11110100_10010010_11111111_11100101_01111101_10111010_10001111_01001000_01011110_01011110_00110011;
assign in[389] = 496'b10011011_10000010_10011011_11101001_11111111_01010101_01110111_01110101_01111000_01110011_10100010_00111110_00000000_11100110_00001001_10111111_00111101_01110011_01101110_11111111_11110011_01011110_00000111_11000111_01111101_01110111_00111010_01101101_00110111_11101011_10111100_01111101_00000100_00011001_10110110_11111100_11111011_00111100_01011101_11111111_11111111_11111111_11111111_10010111_01111101_10000110_11111111_11111111_11111111_10110101_01101111_01000100_11100111_11111111_11111111_10010011_01111000_00111001_11100011_01110110_10001010_11110110;
assign in[390] = 496'b11101011_01110111_11101000_11111111_11111111_11111111_10110010_00111100_11111111_11111111_11111111_11111111_11111111_10000010_00101100_11111111_11111111_11111111_11111111_11111111_00110110_10100100_11000101_10101011_11011100_11111111_11110101_01100110_01101100_01100111_00101011_01011110_11111111_10101011_01111101_00010100_11101100_11110101_01110111_11111001_01001000_00101010_11111111_11111111_10110100_01010001_11111111_00110100_01011110_10001000_10000010_01011110_10111101_11111111_11111011_10101000_10000001_10000010_11010001_11111111_11111111_11111111;
assign in[391] = 496'b01001111_01110010_01111101_01011110_00010001_01101111_10011001_11111010_11110111_11100100_10100101_01000110_00001101_11111111_11111111_11111111_11111111_11111111_01000000_00000011_11111111_11111111_11110010_10100011_11111111_10110110_01011101_11101110_10011111_01001000_01100100_11111111_11111111_00011111_01111101_01111110_01010101_01100011_11111111_11111111_11111110_10110000_10100111_11010011_01100011_11111111_11111111_11111111_11111111_11111111_11011101_01110001_11110111_11100110_10101011_10111000_11110010_11011101_01100011_00110111_01101001_01100000;
assign in[392] = 496'b00010001_11111111_11111111_11111111_11111111_10000111_00010110_11111111_11111111_11111111_11111111_11111111_10101111_00111111_11111111_11111110_11001110_11110101_11111111_11010110_00111111_10101101_01010000_01000010_01011001_11111111_11000001_01110000_00011001_11110000_11111111_00100001_11111111_10101111_01101100_11100111_11111111_11101011_01100000_11111111_10010010_01110101_00001000_11101010_01001010_10010110_11111111_00011110_01101110_00101001_01010110_00000000_11111111_11111111_11110101_10100101_10110010_11111111_11111111_11111111_11111111_11111111;
assign in[393] = 496'b11101001_00011001_01000110_01111001_00110001_11100101_01011101_10000111_10110101_00000011_01010111_11111111_00010110_00000100_11111111_11111111_11111111_11111111_11101110_01100101_11111011_11111111_11111111_11111111_11111111_11001001_00100011_11111111_11111111_11010110_11100100_11111111_11100100_01110111_00100111_00110001_01110101_00000000_11111111_11111111_11001101_10000110_10010111_01011101_10110101_11111111_11111111_11111111_11111111_11010001_01101011_11100101_11111111_11111111_11100000_10100000_00110100_01100001_11111000_01001111_01101010_10011110;
assign in[394] = 496'b11111111_11110100_01111000_11101100_11111111_11111111_11111111_11011011_01010101_11111111_11111111_11111111_11111111_11111111_10101011_00110110_11111111_11111111_11111111_11110101_11001110_00111101_10001011_11111111_11111111_11111111_00011100_00101101_01111100_00111000_01100101_00111011_11111111_11111111_10011010_00101111_11111111_00000101_00010011_11111111_11111110_01010001_10110111_11111111_01010001_11010011_11111111_10110111_00111101_11111111_11111111_00010111_11111110_11111111_00001110_10101010_11111111_11111111_11111111_11110101_11111111_11111111;
assign in[395] = 496'b11111111_10110001_01001010_01111100_00110010_11111111_11001101_01100110_10001110_10111101_01111101_11111111_11011010_01100110_10111001_11111111_10010011_01000101_11111111_00011100_10000001_11111111_11111111_01010000_10001001_11111111_01000101_11011111_11111111_10101111_01100011_11101110_11111111_01001011_11010001_11111111_01010101_10010101_11111111_11111111_00101111_10010100_11001100_01101110_11110001_11111111_11111111_10010111_00101110_01001110_10000100_11111111_11111111_11111111_11011000_01111010_01100010_11110100_11111111_00101011_10010011_11111111;
assign in[396] = 496'b11111111_11010101_01000110_11111111_11111111_11111111_11111111_10011000_00101110_11111111_11111111_11111111_11111111_11111111_10001001_00011000_11111111_11111111_11111111_11111111_11111111_00000010_00001101_11111111_11111111_11111111_11111111_11111111_00011111_10001001_11111111_11111111_11111111_11111111_11111111_00011111_10101100_11111111_11111111_11111111_11111111_11111111_00111110_10110001_11111111_11111111_11111111_11111111_11111111_01000110_10110001_11111111_11111111_11111111_11111111_11111111_00101111_10110001_11111111_11111111_10110111_11011001;
assign in[397] = 496'b11111111_11111111_11111111_11111111_11111111_00001001_00111110_01010000_01000011_10000011_11011010_00100110_10010100_10010111_10100100_10111001_00111100_01101000_11111111_11111111_11010001_01100010_11101111_11111101_00100111_11111111_11111111_11111000_01111001_11100010_11111111_00001101_11111111_11111000_00110101_00100101_11111111_11111111_10100100_01010011_01011101_00011000_11110011_11111111_11111111_00001000_11011101_11101010_11111111_11111111_11111111_11111111_00101100_11111111_11111111_11111111_11111111_11111111_11110110_11111111_11111111_11111111;
assign in[398] = 496'b11111111_11111111_11111111_11111111_11111111_11100101_00100110_01101010_01011110_01101010_10111001_11101100_01011100_10011111_11111101_11111111_10011000_10000010_10100000_00010001_11111111_11111111_11100001_00111101_10010001_10101010_00101010_11111110_11111111_00011010_01111000_11101011_11111100_00100011_01100101_00100110_01111110_00110000_11111111_11111111_11111111_11100000_11000001_01100110_11000011_11111111_11111111_11111111_11111111_10011101_00101001_11111111_11111111_11111111_11111111_11111111_01011001_11010010_11111111_10111101_00110101_11111111;
assign in[399] = 496'b11111111_11111111_11111111_11111111_11111111_00100110_01100100_01100110_01101100_01100110_00011111_01000001_10010101_11110111_11111111_11111111_11101011_01101011_01100000_11111111_11111111_11111111_11111111_00001101_00111110_01011101_10001110_11011001_11010110_00011000_01111011_11001100_11011011_10001010_00011100_00110111_01010110_00010110_11111111_11111111_11111111_11111111_11101001_01011011_11011000_11111111_11111111_11111111_11111111_00001100_00000011_11111111_11111111_11111111_11111111_11000000_01010111_11110110_11111111_01010011_10111101_11111111;
assign in[400] = 496'b00101001_01101100_01100011_01001111_11111111_10100110_01101111_11001110_11110111_01111101_11010011_11111111_00010111_01010111_11111111_11111001_01111101_11010010_11111111_10011010_01101101_11101011_11111001_01101101_11101100_11111111_11011100_01101000_10001010_00011110_01011001_11111111_11110111_11011110_01001000_01111101_01111010_11011001_11111111_00101101_01111101_01111101_01011110_01110111_11001010_11111111_00000001_01111010_10011010_11110100_00111111_01011001_11111111_11111111_00011001_01111101_01111101_01110011_00000100_11000011_10010011_11011111;
assign in[401] = 496'b01010111_00000101_10010011_00101010_11111111_00010100_10011010_11111111_11101001_01011010_11111111_11111111_10101111_00111011_11100010_01000111_10000111_11111111_11111111_11111111_01000110_01111000_10000001_11111111_11111111_11111111_11101111_01011111_01010011_01010010_11101111_11111111_11111111_00110000_10011010_11111111_00001110_00110000_11111111_10100000_00110011_11111111_11111111_11111000_01000001_10101010_10001010_00010101_11111111_11111111_11111010_00101111_10000110_11101110_01001001_01001010_01001000_01011000_00001100_10101000_10110111_11111000;
assign in[402] = 496'b01000100_10110001_10001011_10000111_11111111_00010110_10010101_11111111_11111101_00100001_11111111_11111111_11010101_01010101_11100001_11001011_00011001_11111111_11111111_11111111_10110011_01100111_01100000_11000011_11111111_11111111_11100001_00111010_00010101_01001010_00100000_11111111_11100011_01011001_10101111_11111111_11111000_00100111_10011001_00001010_10010001_11111111_11111111_11111111_10001001_00010110_10001110_00000010_11111111_11111111_11111111_00110111_10011010_11110110_01101000_00001111_11011001_00011100_00101101_10001011_10001111_11001011;
assign in[403] = 496'b00111101_00001110_11111111_11111111_11111111_11010110_01110101_01100100_11100010_11111111_11111111_11111111_11111111_00011000_01111110_10110010_11111111_11111111_11111111_11111111_11010110_01111101_00001110_11111111_11111111_11111111_11111111_11111111_01101101_01100101_11110101_11111111_11111111_11111111_11111111_00101000_01111001_11011110_11111111_11111111_11111111_11111111_00101000_01110111_11101001_11111111_11111111_11111111_11111111_00101000_01111010_11011000_11111111_11111111_11111111_11111111_10001010_01111110_10001000_11111111_11111100_00011000;
assign in[404] = 496'b11111111_11110101_00100111_01110100_10101101_11111111_11111111_00101100_00010111_10111111_10000111_11111111_11111111_11101011_01100000_11111000_10001000_10000111_11111111_11111111_11001001_01011101_11100101_01011000_11011100_11111111_11111111_11101101_01100000_00110011_00001010_11111111_11111111_11111111_11111111_00101110_01110111_11110001_11111111_11111111_11111111_10001010_01011001_01001011_10110111_11111111_11111111_10101101_01011001_10111110_00111001_10000100_11111111_10101010_01000010_11100111_11011011_00010100_11110101_11111111_11111111_11111111;
assign in[405] = 496'b11111111_11101011_10100000_10110101_11101101_11111111_10111011_01110000_01110011_01100000_00100010_11111111_11111111_00110101_01101011_11011000_00011100_01011111_11111111_11111111_00110101_00111111_00111001_01111101_00000101_11111111_11111111_00110101_01111101_01011110_10010100_11111010_11111111_11111111_00000011_01001010_11100011_11111111_11111111_11111111_11111111_11111000_01001100_11100111_11111111_11111111_11010111_11111111_11111111_00110011_11010011_11111111_11111111_00111010_00100101_11110010_00011001_11010011_11111111_01101001_01110001_11100001;
assign in[406] = 496'b11111111_10011111_01100111_01101100_10101010_11111111_10110110_01111011_01101001_11011000_11111111_11111111_11101101_01110010_01111100_11010101_11111111_11111111_11100011_01100011_01111101_01111101_01001100_01001100_00011111_01000110_01111101_01111101_01101100_10000101_00100000_01111101_01111010_01101110_10001001_11101001_11111111_11110011_01101001_01111101_11000001_11111111_11111111_11000000_00111001_01110110_01110101_00100011_00011011_00110110_01111101_01011010_11000011_10000010_00101100_01111010_00101100_10101010_11111011_11111111_11111111_11111111;
assign in[407] = 496'b00000110_00011100_11111111_11111111_11111111_11111111_00000111_00110001_11111111_11111111_11111111_11111111_11111111_00000111_10011011_11111111_11111111_11111111_11111111_11111111_00101100_00001011_10100100_00011010_00110110_11111111_11111111_01011111_10101110_10110010_10110010_01010000_11111111_11100000_01110101_11110001_11111111_11111001_01100011_11111111_10101101_00110001_11111111_11111111_10101101_00110100_11111111_01000100_10101001_11111111_11111111_10001001_10001011_11000010_01001001_11110001_11111111_11111111_10111001_11111111_11111111_11111111;
assign in[408] = 496'b11111111_00110111_10101100_11111111_11111111_11111111_10101101_01111110_00011111_11111111_11111111_11111111_11111111_11000111_01001111_00011111_11111111_11111111_11111111_11111111_11111111_01001101_00001110_11111111_11111111_11111111_11111111_11111111_01001101_10010101_11111111_11111111_11111111_11111111_11111111_01001101_10010101_11111111_11111111_11111111_11111111_11111111_01001101_10010101_11111111_11111111_11111111_11111111_11111111_01100011_10010101_11111111_11111111_11111111_11111111_11111111_01101001_10010101_11111111_11111111_00101101_10010101;
assign in[409] = 496'b11111111_11111111_11111111_00000110_01110001_11111111_11111111_11111111_10111011_01111100_10011001_11111111_11111111_11111111_11100111_01101000_00011001_11111101_11111111_11111111_11111010_00111110_01000101_11111111_11111111_11111111_11111111_00000100_01101010_11011000_11111111_11111111_11111111_10111001_01110111_10101000_11111111_11111111_11111111_11100111_01100100_00100110_11111111_11111111_11111111_11111111_00001001_01010001_11010001_10000111_01101010_01111100_00001101_01100010_01111101_01110001_00100101_10011001_10011111_11111111_11111111_11111111;
assign in[410] = 496'b10101001_01100100_01111101_01011001_10101011_11101110_01011101_00101111_10111001_00000000_01110000_11111111_11110100_01101011_10000010_11111111_11111110_00110001_11111111_11111111_00011101_01100011_11011000_00110010_01010101_11111111_11111111_10110000_01111101_01101110_00110110_11100111_11111111_10110011_01010010_01111101_00110010_11111111_11111111_00001001_01111000_00111001_10011001_01100000_11111111_11111111_01110000_10011101_11111111_11100100_01101010_11111111_11111111_10111101_11011100_11111010_00010001_00110101_11111111_01100110_01010000_11011110;
assign in[411] = 496'b00100101_10011101_00100000_01000100_11100011_10011010_11111111_11111111_11111111_10010000_10010100_00010001_11011110_11111111_11111111_11111111_10101011_10011100_10001001_11000101_11111111_11111111_11111011_00110001_11011000_11101111_00110101_10000011_00010101_01001000_10000100_11111111_11111110_01000001_10001110_10110111_10100111_01010011_10111110_11110101_01000010_11111111_11010010_11111100_10110011_00110001_11111110_00011100_10001001_01100000_11110100_00110111_10111001_11111111_11111111_10101011_00001110_00100110_00000001_11110111_10000100_10110111;
assign in[412] = 496'b11111111_11111111_11111111_11111111_01010001_11111111_11111111_11111111_11111111_10010010_01111011_11111111_11111111_11111111_11111111_10111010_01110100_01000101_11111111_11111111_11111111_11001111_01011011_01100010_11101010_11111111_11111111_11101010_01011011_01110010_11001101_11111111_11111111_11111110_00101110_01111100_10010101_11111111_11111111_11111111_10010000_01111101_00000101_11111111_11111111_11111111_11010000_01110001_00100000_11111111_11111111_11111111_11111111_00011101_01100000_11111010_11111111_11111111_11111111_11111111_11111111_11111111;
assign in[413] = 496'b11111111_11111111_11111111_11111111_11111111_11111111_11110100_10111000_00011010_00011010_00011010_11111010_00110101_01111010_01111110_01111101_01111101_01101110_01001001_01111101_00011001_10111111_11110010_11110010_11110110_01111000_10010011_11111110_11111111_11111111_11111111_10000011_01110011_11011101_10010011_11101001_11111111_10100101_01101101_01111011_00111010_01001100_11110001_10001110_01101001_00101100_01111101_01111110_01010000_00100010_01111101_00100000_11100100_10101100_10001100_01100001_00111010_10110111_11111111_11111111_11111111_11111111;
assign in[414] = 496'b10010010_01011101_10010001_11111111_11111111_10101001_01001101_11010001_01001101_10001111_11111111_11111100_01000110_11011110_11111111_11101110_01011100_11110101_11000000_00100001_11111111_11111111_11111111_00111010_10100111_10010101_10011110_11111111_11111111_11111111_00011010_10000010_10111010_10011101_11111111_11111111_11111111_00011010_10000001_11101010_00011111_11111111_11111111_11111111_01001010_11000000_11111111_00110010_11111101_11111111_11000000_01011000_11111111_11111111_10011000_10001000_11111100_00111110_00010100_00001110_00111010_00101001;
assign in[415] = 496'b11111111_11111111_11111111_11111111_11111111_11111110_00011010_01111101_01010101_00111111_10000111_11100011_01001101_01110111_01110110_01111101_01001001_01111001_01001101_00100011_11011011_00111111_01011001_11101110_01010001_01111101_00011110_01101001_00100111_11101010_10111101_01111101_01000011_01011010_10101101_11111111_11111111_00000011_01110001_11111111_11111111_11111111_11111111_11000110_01101110_00101000_11111111_11111111_11111111_10111111_01011000_00100001_11101111_11111111_11111111_10100100_01110110_00000111_11111111_01111011_00010111_11111111;
assign in[416] = 496'b11111111_11000000_00011010_01101001_01111101_11101010_00100000_01110100_01111101_01000111_00010111_11110110_01000111_00110011_11011100_11000100_11111111_11111111_00000000_01010010_11101100_11111111_11111111_11111111_11111111_00110111_00001101_11101101_10101010_00100000_00011101_11111111_00011100_01011010_01101101_01111101_01111011_01001000_11111101_10001001_01110001_00010111_10100010_11100000_11111111_11111111_01110110_10110010_11111111_11101000_11110110_11111111_11111111_01110111_00000011_00111100_01111000_10110010_11111111_01001001_10001011_11110110;
assign in[417] = 496'b11111111_11111111_10011011_01111000_11001100_11111111_11111111_11011001_01110111_00000110_11111111_11111111_11111111_11011011_01011100_01110000_10100001_11101010_11111100_00100110_01111001_01101010_01100100_01110100_01101010_11111111_10001000_01101110_11100001_11111100_10110100_01111101_11100011_01110010_10010110_11111111_11110110_01001010_01000100_00101011_00111101_11111001_11111111_00101100_01010000_11100010_01110101_11100001_11111111_11100110_01010011_11100001_11111111_00010011_11111111_11111111_11111111_11111001_11111111_11111111_11111111_11111111;
assign in[418] = 496'b11100101_00001010_01101110_01101011_00101101_11010100_01101000_01010011_00100100_01001000_01111110_11010100_01100110_00010110_11111110_11111111_11111100_01101010_01010010_00101111_11111111_11111111_11111111_11111111_01001001_01101111_11101100_11111111_11111111_11111111_11111111_01000100_01100100_11110110_11111111_11111111_11111111_11010101_01110111_01111011_00000001_11111101_11100101_11011110_00011011_00000000_00000000_01111110_01000000_00100100_01110100_01101000_11001011_11111110_10101100_01010111_01111110_01110111_10101110_00100010_01100010_10101111;
assign in[419] = 496'b11111111_11111111_11110101_00110110_01111101_11111111_11111111_11111111_11001100_01111101_01111100_11111111_11111111_11111111_11101000_01010010_01111011_10011011_11111111_11111111_11111011_00111001_01111010_10001010_11111111_11111111_11111111_10000001_01111101_00011100_11111111_11111111_11111111_10111101_01111010_01001110_11110010_11111111_11111111_11111101_01010100_01110010_11010010_11111111_11111111_11111111_10101000_01111101_00001110_11111111_11111111_11111111_11111111_00110011_01110011_11101111_11111111_11111111_11111111_11110101_11111111_11111111;
assign in[420] = 496'b11111111_11111111_11110001_01010001_01100000_11111111_11111111_11111101_00110110_01110100_11011111_11111111_11111111_11111111_00011101_01110011_10111100_11111111_11111111_11111111_10101010_01111010_10110100_11111111_11111111_11111111_11001010_01110010_00100000_11111111_11111111_11111111_11011111_01100000_01010100_11101111_11111111_10111110_10010111_01010101_01101011_10001001_10010010_01001110_01111101_01111100_01111101_01111100_01111100_01111101_00110001_10101101_11010101_10101011_11001010_10011100_11001100_11111110_11111111_11111111_11111111_11111111;
assign in[421] = 496'b00010000_10010001_10111100_10010010_10110111_11001110_00100100_11111111_11111111_11111111_11111100_11111111_10001101_10110010_11111111_11111111_11111111_11111111_11111111_10110110_10011000_11111111_11111111_11111111_11111111_11111111_11100110_00101010_11111111_11111111_11111111_11111111_11111111_11111111_00001011_00111100_01000101_10001011_11111111_11111111_11111111_11111111_11111001_10000110_00001001_11111111_11111111_11111111_11111111_11111111_10010101_00001001_11111111_11111111_11111111_11101000_00000000_00010010_00001001_11111111_11011101_10000011;
assign in[422] = 496'b11000011_10100001_11000011_11111110_11111111_01010101_01100100_01000011_01111100_01010101_11011001_01010100_10010101_11110011_11100101_01000111_01110101_01001001_01000111_11111111_11111111_11111111_00010100_00000111_01011111_01010011_11111010_11111111_11100000_01110101_11011011_00000110_01001100_01011111_00111011_01110101_10011010_11111111_00110010_11111010_10100011_10001110_11001000_11111111_11100101_01110110_11111111_11111111_11111111_11111111_11111111_00101111_00111101_11111111_11111111_11111111_11111111_10101000_01101011_10100101_00100010_01101000;
assign in[423] = 496'b11111111_11111111_11111111_10100011_10000110_11111111_11111111_11111111_11111110_00101110_11000110_11111111_11111111_11111111_11111111_10100000_00101100_11111111_11111111_11111111_11111111_11101110_01011101_11001010_11111111_11111111_11111111_11111101_00110001_00010000_11111111_11111111_11111111_11111111_10100100_01100110_11110000_11111111_11111111_11111111_11100111_01100110_10111011_11111111_11111111_11111111_11111111_00101001_00011101_11111111_11111111_11111111_11111111_10101000_01000001_11110101_11111111_11111111_11111111_11111111_11111111_11111111;
assign in[424] = 496'b11111111_11010101_01111101_10101011_11111111_11111111_11111111_11101111_01111110_10100101_11111111_11111111_11111111_11111111_11101111_01111101_10100110_11111111_11111111_11111111_11111111_11001011_01111110_11011110_11111111_11111111_11111111_11111111_10100111_01001011_11111111_11111111_11111111_11111111_11111111_00110111_00100011_11111111_11111111_11111111_11111111_11011110_01110110_10000111_11111111_11111111_11111111_11111111_11001010_01110100_11100101_11111111_11111111_11111111_11011011_00110101_00110111_11111111_11111111_10000001_11101000_11111111;
assign in[425] = 496'b11111111_11111010_00110011_01011101_11111001_11111111_11111111_11111111_01010000_10011100_11111111_11111111_11111111_11111111_10011100_00111011_11111010_11111111_11111111_11111111_11101101_01101100_11010000_11111111_11111111_11111111_11111111_00010101_10001000_11111111_11111111_11111111_11111111_11101011_01101100_11110110_11111111_11111111_11111111_11111111_10000011_00001011_11111111_11111111_11111111_11111111_11111001_01010100_11000001_11010110_10001001_11010101_11111111_11111010_00100111_01010111_00111000_10001101_11100001_11111111_11111111_11111111;
assign in[426] = 496'b11111111_00001110_01101010_11111001_11111111_11111111_11110010_01100011_11000000_11111111_11111111_11111111_11111111_00001110_01000111_11100100_11111111_11011101_11001111_01011100_01111111_01011100_01101010_01000111_01100011_11111111_01100011_10001111_11111111_11110010_01100011_01011100_11001000_01011100_11111111_11111111_00000111_00111000_11111111_00100011_10001000_11111111_11110010_01110001_11101011_11111111_01111000_11111001_11111111_10001111_00011100_11111111_11111111_00001110_11111111_11111111_11010110_11101011_11111111_11111111_11111111_11111111;
assign in[427] = 496'b11111111_11111111_11111111_11111111_11111111_11111111_11000000_01001101_01101111_01111101_00110100_11111111_10011010_01011101_00000100_00101010_01011100_01101100_11011000_01001100_11110001_11000111_01101110_00101100_00101110_11000001_01011001_10001111_01100001_10110001_01101000_10101111_11111111_10010101_10001010_11101100_00100011_00111110_11111010_11111111_11111111_11111111_10001000_01101001_11101000_11111111_11111111_11111111_10111110_01101110_11001100_11111111_11111111_11111111_11011001_01011011_11000000_11111111_11111111_10110010_11111111_11111111;
assign in[428] = 496'b10010001_01111100_00001001_11111111_11111111_11111111_11010000_01110101_01110100_11000100_11111111_11111111_11111111_11111111_00001011_01111100_00100011_11111111_11111111_11111111_11111111_10000011_01111011_00100010_11111111_11111111_11111111_11111111_00111111_01111100_00000010_11111111_11111111_11111111_11001011_01111100_01110110_11001101_11111111_11111111_11111111_10111000_01111100_01101010_11111111_11111111_11111111_11111111_00010000_01111101_00111110_11111111_11111111_11111111_11111011_01010111_01100001_10101101_11111111_00110110_11110110_11111111;
assign in[429] = 496'b11100101_11111111_11111111_11111111_11111111_11111111_01010100_11101010_11111111_11010100_00011100_11111111_11111100_01101000_11101010_10001001_01100000_10100111_11111111_11111110_01011010_01011011_00100111_11110110_11110011_11111111_11110110_01011001_01101011_00000101_00111110_00110101_11110001_00111101_00011000_11011001_10111000_11010111_11111110_00000010_01000101_11101111_11101111_11111111_11111111_11111111_01101100_01001000_01101000_01100101_11111101_11111111_11111111_01011111_00011001_01101110_10011000_11111111_11111111_11110010_11111111_11111111;
assign in[430] = 496'b11111111_11100010_01100111_01010111_11101111_11111111_11011001_01011110_01011001_11100110_11111111_11111111_11111100_01010010_01010111_11100101_11111111_11111111_11111111_00010110_01110000_11001110_11111010_10110011_10010000_11001111_01111100_00001011_00000001_01100010_01011010_01101010_00110111_01111101_01111100_00100110_11000110_11110111_01001100_01111101_01111101_10011001_11111111_11100011_01000110_00011001_01111101_00110101_11110011_10000001_01100100_10010111_11111111_00110110_01001000_01011111_00010110_11100000_11111111_11111111_11111111_11111111;
assign in[431] = 496'b10001101_01010111_01110010_01011000_01111010_10101011_00011110_11011000_11110110_11100011_00001101_11111111_01100000_10010001_11111111_11011001_00110111_01010100_11111111_00100000_00110000_10101011_01100100_00011101_11101111_11111111_00001010_01111000_01011011_11010011_11111111_11111111_11010011_01110001_01110011_00011110_11111111_11111111_11111111_00111000_10100010_10100011_01111100_10011001_11111111_11111111_01001011_01010010_00000101_01010011_01110100_00011101_11110101_10101001_01110100_01111101_01111110_01111101_01101011_11010010_10101001_10000001;
assign in[432] = 496'b11111111_11111111_11111111_11111111_11111111_11111111_11010011_00100101_00110111_00011111_11000110_11111011_00011010_01011100_00010000_01111101_10000110_01110001_10010001_01100000_11000101_00101000_00011010_11111010_01110101_11011101_01000000_00101111_10101000_11111100_10100101_01001101_11111111_11111111_11111111_11111111_11011000_01100011_10111010_11111111_11111111_11111111_11001000_01101111_10101111_11111111_11111111_11111111_11010100_01101110_10110101_11111111_11111111_11111111_11101000_01100000_10011000_11111111_11111111_10101000_11111111_11111111;
assign in[433] = 496'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11010101_00001001_01100000_10001100_10010000_10111010_00000101_01110010_00010100_10011101_10111010_10100111_01110111_01101111_01101111_00111000_01101011_11111111_10011111_00011101_11111101_11101100_11000100_11011010_11111111_00111000_11101101_11111111_11111111_11111111_11111111_11111000_01011111_11111111_11111111_11111111_11111111_11111111_11111111_00101011_11010001_11111111_11111111_11111111_11111111_11111111_11011101_01001001_10010000_10111100_11100111_11110101_10100110_00010100;
assign in[434] = 496'b01000101_01101101_01010000_00101001_10001110_01110101_10100101_11011101_11011101_10110110_01100101_00011110_01111101_11001001_11111111_11111111_10110100_01100111_11010001_01110101_01101010_11001001_00010010_01111001_00000110_11111111_11001010_01101101_01111110_01111101_10101101_11111111_11111111_00010100_01111000_01000000_01111100_00100001_11101001_00000101_01101110_10111111_11111111_10101100_01101110_01001101_01100011_11000100_11111111_11111111_11111111_11011011_01100011_11110001_11111111_11001001_11000001_10000011_01010100_01110010_01100001_00010101;
assign in[435] = 496'b11111111_10100111_00111111_01110010_01010001_11111111_11101001_01110011_10100111_11111001_10000111_11110110_11111111_11101001_01111110_11100110_11011100_01011101_11111111_11111111_11111111_01000011_01000110_01011001_10011110_11111111_11111111_11101010_01001001_01111110_10100110_11111111_11111111_11011110_01011011_00001101_01010100_10101011_11111111_10111100_01100111_10011101_11111111_00111010_10101001_11111111_01101111_10111110_11111111_11101000_01011111_11101010_11111111_00000111_11100111_11011011_01000100_10100110_11111111_00110011_11100011_11111111;
assign in[436] = 496'b10011000_01111010_10101011_11111111_11111111_11111111_01100011_01111011_10000001_11111111_11111111_11111111_11111111_01100010_01111010_00010010_11111111_11111111_11111111_11111111_00111010_01111011_01100100_11111111_11111111_11111111_11111111_10000011_01111010_01100011_11111111_11111111_11111111_11111111_10000011_01111011_01101110_11100010_11111111_11111111_11111111_11101000_01111010_01100011_11111111_11111111_11111111_11111111_11101000_01111011_01111000_11000011_11111111_11111111_11111111_11111111_00101111_01100011_11111111_11111111_11011101_10000001;
assign in[437] = 496'b11111111_11111111_11011111_01011001_01100001_11111111_11111111_11111111_11111111_10000011_01110111_11111111_11111111_11111111_11111111_10101010_01111101_10100011_11111111_11111111_11111111_11100011_01101111_00011010_11111111_11111111_11111111_11111111_00110100_01011101_11110110_11111111_11111111_11111111_10010000_01110010_11001111_11111111_11111111_11111111_11100000_01010010_00001011_11111111_11111111_11111111_11111100_00111011_01000111_11101110_11111111_11111111_11111111_10001010_01110001_11100101_11111111_11111111_11111111_11111111_11111111_11111111;
assign in[438] = 496'b11111111_11100000_01011001_01100011_11001010_11111111_11111111_10010110_01111011_01111100_10111011_11111111_11111111_11111111_00001101_01111100_01010110_11111111_11111111_11111111_11101111_01100111_01111011_00011010_11111111_11111111_11111111_10010111_01111101_01111100_10100001_11111111_11111111_11111011_00111011_01111100_01100100_11110110_11111111_11111111_11001111_01111011_01111100_00000010_11111111_11111111_11111111_10010011_01111100_01100110_11100001_11111111_11111111_11111111_01110001_01111011_00001001_11111111_11111111_01011010_11000010_11111111;
assign in[439] = 496'b11101001_00100000_01101100_01010001_10011101_11001100_01101001_01001100_10010001_10000010_01100011_11101010_01011001_00011001_11101010_11111111_11111111_11100011_10101010_01111010_11110111_11111111_11111111_11111111_11111111_11011101_01010101_10001111_11011010_11111111_11111011_11110100_11111111_11100110_00111100_01111000_00111110_01010011_01000101_11111111_11111111_11111111_00110000_01110001_00010110_11001011_11111111_11111111_00001001_01110100_10111100_11111111_11111111_11111111_11111101_01101101_01000011_11000000_10111011_11010101_00100110_01111110;
assign in[440] = 496'b11111111_10011101_01111011_01111100_01111011_11111111_11111111_10111111_01111100_01100101_01111100_11111111_11111111_11111111_11110001_01111011_01111100_01111011_11111111_11111001_11001001_00001111_01111011_01111100_00100001_11101001_00010011_01111101_01111010_01100010_01111101_00010010_01001111_01111011_01101001_10011000_11010000_01100010_00011011_01101111_10101011_11011100_11111111_11001011_01111010_00001101_01111100_01111011_01111100_01000110_01101000_01111100_10101111_01000110_01111011_01111100_01111011_01101110_00100111_10000110_10000110_11100101;
assign in[441] = 496'b11111111_11100110_00010111_01011000_00101010_11111111_10001100_00111110_11000001_10011101_11100001_11111111_00010011_00000101_11111111_11111111_11111111_11111111_11100010_01000000_11111111_11111111_11111111_11111111_11111111_11111111_00010101_00110000_10001011_10001101_10011110_11011010_11111111_11111111_11011011_10110011_01000011_00101101_11101001_11111111_11111111_11111111_10101111_00011100_11111111_11111111_11111110_10100000_00111101_01100110_11011011_11111111_11111111_10111100_00000000_10011110_10011011_11111111_11111111_10000011_11001110_11111111;
assign in[442] = 496'b10010100_00110100_01000100_01111100_01011000_00111100_01111110_01111101_01010100_01111101_01101101_10010111_01111100_00110111_11111011_11111111_11111111_11111111_11010000_01111000_00111000_11111011_11111111_11111111_11111111_11111111_10000111_01111101_01100010_10010100_11101001_11111111_11111111_11111110_10010011_01111000_01111110_01101011_10111000_11111111_11111111_11111111_11111011_10011001_01111010_01011101_11111111_11111111_11111111_11111111_10111110_01111010_01011110_11001101_10101110_10010100_00110100_01111101_01110101_01011001_01111101_00110101;
assign in[443] = 496'b11111111_11111111_11111001_00000001_10011110_11111111_11111111_11111111_11000101_01111100_01111100_11111111_11111111_11111111_11111111_11110001_01100101_01111100_11111111_11101001_10111100_00010010_01000010_01111010_01111100_00101100_01111010_01011100_00111000_10000010_00101111_01011010_01001110_11000100_11111110_11111111_11111111_00001011_00100010_00101111_11101111_11111111_10111110_11001111_01000011_01001101_10111000_11111111_10111000_01101011_01111100_01111100_11000100_11111111_11111111_11111111_11010000_10001001_11001001_11111111_11111111_11111111;
assign in[444] = 496'b01111011_01111110_01111011_00010010_11101000_01111101_01010101_01000011_01111000_01111101_01010001_01111101_00110100_11111001_11111111_11110011_10011001_01110000_01101100_11101100_11111111_11111111_11111111_11111111_00110101_01011001_11111111_11111111_11111111_11111111_11111111_00001101_01101000_11110001_11111111_11111111_11111111_11111111_00010110_01111101_10100010_11111011_11110100_11111111_11111000_01100001_01100010_01100110_01010111_00011000_11110010_00011111_01111010_11011011_01000110_01111100_01111110_01111101_01111101_11000000_01011001_01111100;
assign in[445] = 496'b01100100_00100010_10001111_10100001_11110101_10010100_11100100_11111111_11111111_11111111_11111111_01110110_10111000_11111111_11111111_11111111_11111111_11111111_10000011_01011010_10111011_11001101_11111111_11111111_11111111_11111100_10011010_01010000_01110110_01010000_10000100_11100001_11111111_11111111_11111111_11100101_10010100_01011001_00111010_11111111_11111111_11111111_11111111_11111111_11001011_01111101_11111111_11111111_11111111_11111111_11111111_11000111_01111100_11111111_11111111_11111010_01010001_01100111_01111011_11111111_11101101_10011110;
assign in[446] = 496'b01110001_11011101_11111111_11111111_11111111_01100011_10001111_11111111_11111111_11111111_11111111_10100100_01101010_11111001_11111111_11111111_11111111_11111111_11000000_01000111_10001000_01010101_01010101_00110001_11100100_11000000_01111111_00001110_10101011_10001111_00110001_01100011_00011100_00010101_11111111_11111111_11111111_10100100_01111111_01000111_10101011_11111111_11111111_11111111_10010110_01111111_00111000_00011100_11001110_10001000_01001110_01111111_00011100_11010110_01000111_01110001_00111000_00001110_11001111_11111111_11111111_11111111;
assign in[447] = 496'b11111101_11110001_11110001_11110001_11110100_10100001_01000010_01111100_01111011_01111011_01110001_01100010_01111101_01110001_01001111_01001110_01001110_01100110_01111011_00010011_11101000_11111111_11111111_11111111_11100010_01010000_11101110_11111111_11111111_11111111_11111111_11111111_00001110_11111111_11111111_11111111_11111111_11111111_10101111_00010111_11111111_11111111_11111111_11111111_11101001_01110000_01101101_10110100_10000011_00111010_11011011_01010011_01111101_01000101_01111100_01111011_10010010_11111010_00110001_11100110_11111111_11111111;
assign in[448] = 496'b11111111_11111110_10000111_01100111_01111101_00010010_10011010_00110001_01111101_01111101_01111101_10010000_01100101_01111101_01111101_01111100_01110101_01011100_11111111_10010110_01111101_01001011_11001001_11011011_11111111_11111111_00111110_01110001_10111000_11111111_11111111_11111111_11111111_01101001_00000110_11111111_11111111_11111111_11111111_11001011_01111011_10001111_11111111_11111111_11111111_11111111_11111010_01010110_01011101_10111001_11111111_11111111_11010110_11111111_10101111_01100010_01110111_00110101_00100001_11111011_00001111_01100101;
assign in[449] = 496'b10111011_00011000_01000101_01000110_01000101_01001001_01111100_01111101_01111100_01111101_01111100_01111100_01111011_01000000_10100110_10101100_11100000_01111011_01111100_10001101_11111000_11111111_11101101_11111111_10011011_01110001_11111111_11111111_11111111_11011000_11000010_10010110_00101000_11111111_11111111_11101011_00101001_00110101_01101000_01111101_10100110_10100110_01001100_01111100_01111101_01111100_01111100_01111011_01111011_01111100_01111011_01111100_01111011_00001101_01000110_00110011_11000000_00010110_01111100_11111111_11111111_11110001;
assign in[450] = 496'b11110000_01100000_01111111_10110000_11111111_11111111_00100000_01111111_01000000_11111111_11111111_11111111_11000000_01111111_01101111_11010001_11111111_11111111_11111111_00101111_01111111_00010000_11111111_11111111_11111111_11010000_01111111_01111111_11110000_11111111_11111111_11111111_00000000_01111111_10010001_11111111_11111111_11111111_11111111_01101111_01111111_00100000_00000000_01000000_01000000_01100000_01111111_01111111_01111111_01111111_01111111_01111111_01000000_10100000_00000000_10010001_11010000_11100000_11111111_11111111_11111111_11111111;
assign in[451] = 496'b11010001_01100100_01000001_00011101_00111100_11000001_01100100_11000110_11111111_11111111_11111111_11111111_01001011_10001011_11111111_11111111_11111111_11111111_11101010_01101111_11101110_11000001_00100111_00110001_11111110_11110100_01011111_01010000_01100000_00100000_01110001_11110011_11111111_11010000_10011011_11111001_10110101_01010101_11111111_11111111_11111111_11111111_11111111_10011011_00011000_11111111_11111111_11111111_11111111_11011011_01000011_10011011_11111111_10000010_10000010_00011000_01110100_01000110_10111011_10000001_11010101_11111111;
assign in[452] = 496'b11111111_11000011_01111101_01111101_01111101_11111111_11111111_11111001_01000100_01110100_01000001_11111111_11111111_11111010_11011111_01011010_01111101_01111101_11101010_10001011_01011100_01111101_01111101_01111101_01110101_01101101_01111101_01100010_00010111_11010011_01011000_01001000_01100100_00001110_11100101_11111111_11111100_01001111_00011000_00010010_00011110_00111000_10011100_00101110_01111010_10101011_01111101_01111101_01111101_01111101_01111101_01010001_11100100_10000111_10000010_00101010_01111110_01100100_10111000_11111111_11111111_11111111;
assign in[453] = 496'b01111001_01100110_01001110_00011101_11111111_01111010_01010110_11100110_11111111_11111111_11111111_11000101_01111100_10001010_11111111_11111111_11111111_11111111_11110010_01010101_01101101_11001001_11111110_11111111_11111111_11111111_11100111_01000100_01111110_01010010_00111000_11001110_11111111_11111111_11111011_00010001_01111100_01110110_10101110_11111111_11111111_11100010_01100011_01101010_10110000_11111111_11111111_11111111_00000010_01111101_01000111_01010110_10000110_11111111_11111111_10101101_01111011_01111100_01101001_11111111_11010010_10110010;
assign in[454] = 496'b10010010_01011001_01111101_01111101_00010110_01110111_01111101_01100000_01000010_01001011_01111101_01100101_01111010_10010010_11111001_11111111_11011011_01111101_01111101_00111011_11111111_11111111_11111111_10111000_01111101_01111110_10000111_11111111_11111111_11111110_01000110_01111110_01111101_00001111_11111111_11111111_11010010_01111101_01110110_01111101_00111011_11111111_11100011_01011111_01111101_00111011_00100100_00111110_10100111_01100111_01111101_01110000_11001001_10110100_01111101_01101100_01111110_01101111_10001111_01110110_11000011_11101100;
assign in[455] = 496'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111001_10011100_11011011_11110111_11111111_11000010_00010100_01100100_01101100_01111101_01101001_01100000_01111101_01111101_01111101_11110101_01000101_01111101_01111101_01000111_01000111_00100001_11000110_01111101_01111101_11001001_11111111_11111111_11111111_11100010_01111101_10000100_11111111_11111111_11111111_11111111_11101101_01110011_00110100_10100110_10110100_11010100_11111111_11111111_10100110_01101100_01111110_01111101_01011001_11110100_11010000_10110010;
assign in[456] = 496'b11111111_11111111_11001110_10101110_11100111_11111111_11111111_11111111_01000000_01011000_01010011_11111111_11111111_11111111_11111111_01000110_11000110_00110000_11111111_11111111_11111111_11111111_00001001_00111101_01101000_11010110_10101110_10101011_10011110_10011110_01101000_00110111_01100011_00111011_00110111_01010001_01000110_01111010_10010100_11111111_11111111_11111111_11100010_10001011_01111000_11010001_11111111_11111111_00011011_01111010_01111101_01000010_11111111_11111111_11111111_11110000_10100001_11000000_11110100_11111111_11111111_11111111;
assign in[457] = 496'b11111111_11111111_11111111_11111111_11111111_00110100_01111100_01111101_01010011_11001000_11111111_01110010_01111110_01111101_01111110_01111101_01110010_10101101_01111100_01111101_01100011_10011001_11010111_01101101_01000100_10101000_10101000_11101011_11111111_11111111_01011000_01011001_11111111_11111111_11111111_11111111_11111011_01011101_01011001_11111111_11111111_11111111_11111111_11100111_01110010_01000101_11111111_11111111_11111111_11111111_10010101_01111100_10101101_11111111_11111111_11111111_10101110_01111100_01010100_10111110_01111101_01111100;
assign in[458] = 496'b10010010_10000010_10000010_10000010_11001110_01010111_01111101_01111101_01111101_01111101_01111101_01110110_01111101_01110100_10000100_10111110_10101010_01111101_01111101_01111101_01011001_11100110_11111111_11111011_01101110_01111101_01011011_11011010_11111111_11111111_10101001_01111101_11001101_11111110_11111111_11111111_10111110_01110100_01111101_11111111_11111111_11111111_11100111_01101001_01111101_01011111_11111111_11111110_10011101_01110010_01111101_00100010_11100000_11111111_00000010_01111101_01111101_01011100_11110010_01111101_01011111_11010011;
assign in[459] = 496'b11010010_01010000_01110101_01000000_01100010_11101101_01010111_00111011_11110111_11111111_11001100_11111111_00110001_01010000_11110111_11111111_11111111_11111111_11101111_01110011_10100111_11111111_11111111_11111111_11111111_11110111_01101111_11010001_11111100_10111011_01010000_10111100_11111111_00011100_01000101_01100100_01111100_00111010_11101110_11111111_11111111_11011011_01011010_00101110_11111110_11111111_11111111_11111111_10100101_01111101_00010110_10100010_11001000_11111111_11110101_01101100_01110110_01100100_01001100_10010101_11011011_11111100;
assign in[460] = 496'b11111111_11111101_11111001_11111001_11111001_11001110_00100001_01010111_01111101_01111101_01111101_10001010_01111101_01111101_01111101_01111101_01110000_01110011_01111101_01111010_00111000_10011100_00000100_11001101_00010011_01111101_00100100_11111111_11111111_00001111_00111000_01101001_01111101_00010100_11111111_10100100_01110111_01111101_01111101_01111101_10000010_10011000_01110111_01111101_01111101_01001000_01111101_01110101_01111101_01010001_00010101_00010000_11101110_00111001_01111101_01011101_10111101_11111111_11111111_11111100_11111111_11111111;
assign in[461] = 496'b11111111_10011001_01111100_11001011_11111111_11111111_11111111_01100000_01000000_11111010_11111111_11111111_11111111_10101010_01111100_10011001_11111111_11111111_11111111_11110110_01011110_01001110_11111110_11111001_11111001_11111111_10000110_01111100_01110010_01110001_01110001_01110110_11001111_01110111_00011011_11111111_11111111_11111111_11000110_01001111_01001100_11110001_11111111_11111111_11110101_00101101_01110111_11001110_11111111_11111111_11111111_10000111_01110101_11001001_11111111_11111111_11111111_11111111_10001010_11111111_11111111_11111111;
assign in[462] = 496'b11001100_01110111_01010000_11111011_11111111_11111111_10011011_01111100_10100011_11111111_11111111_11111111_11001010_01111000_00100011_11111111_11111111_11111111_11111101_00111010_01111110_11010101_11111111_11111111_11111111_10011011_01111001_01111110_01010100_01000001_01010000_01011111_01011111_01110000_00000001_10100001_10101001_00011010_01111110_01111111_10011010_11111111_11111111_11101111_01000000_01011011_00001010_11111110_11111111_11111111_00101101_01110100_11001101_11110000_11111111_11111111_11111000_00111011_10101001_11111111_11111111_11111111;
assign in[463] = 496'b11111111_11111111_11111111_11111111_11111111_10001010_00110100_01110010_01111100_00010101_11001101_01010011_01111110_01111101_01111110_01111101_01111101_01111000_01111100_01111101_01111100_01110011_11010111_10001111_01111100_01111101_01111110_01111101_00001100_11111111_10111000_01111101_01111100_01101001_10000100_11111111_11111111_10000101_01111100_11011100_11110001_11111111_11111111_11111111_00010000_01111101_11111111_11111111_11111111_11111111_11011101_01010011_01110111_11111111_11111111_11111111_11101100_01001001_01111100_11111111_00010000_01111100;
assign in[464] = 496'b11111111_11111111_11111111_11111111_11111111_00000100_01100111_01110000_01000101_11011010_11111111_01000111_10111000_11111111_11111111_11000011_01001111_11000111_11010000_11111111_11111111_11111111_11111111_10101101_10010000_11101101_11111111_11111111_11111111_11110001_00001001_00100011_00101111_00000010_10010011_00001010_00111010_00010100_00000101_11101000_11010110_11110011_11111111_11111111_10011011_10101111_11111111_11111111_11111111_11111111_11111111_00110100_10110100_11111111_11111111_11111111_11111111_11111111_01001011_11111111_11111111_11101100;
assign in[465] = 496'b11111111_11111100_10001000_01111110_01010101_11111111_11111111_11100011_01111010_00111110_01000111_11111111_11111111_11111111_10010011_01111110_01001010_01110111_11111111_11101000_10011110_01101101_01111110_01000001_11101001_11000111_01100100_01111111_01001000_00010010_00111010_11111111_01111100_01010110_10110101_11111101_10101001_01101111_11110110_00111011_11101110_11111111_11111111_10101000_01110111_11101011_00110010_10001000_10001010_10111011_00100000_01101100_11110110_01011100_01001100_01101000_01111110_01111110_00000010_11111011_11010011_10111100;
assign in[466] = 496'b11111111_11111111_11111111_11111111_11111111_00001111_01001101_01111101_01111100_01010110_11010110_01000101_01111100_01111100_01111101_01100000_01110111_01011001_01111110_01111101_01111101_01110001_11100101_00001101_01111101_10100100_01100001_01011101_10011011_11101110_01011111_01111000_11111111_11111111_11111111_11111111_10011110_01111110_00000101_11111111_11111111_11111111_11101000_01100001_01111101_11000110_11111111_11111111_11111111_10000011_01111100_00010100_11111111_11111111_11111111_11100011_01111110_01100000_11001000_01000101_01111101_10001001;
assign in[467] = 496'b11111111_11111111_11101010_01011100_00010000_11111111_11111111_11111101_00011100_01110111_10100100_11111111_11111111_11111111_11001000_01111101_00011000_11111111_11111111_11111111_11111111_00111010_01110111_11100100_11111111_11111111_11111111_11111001_01110010_00001011_11111111_11111111_11111111_11111111_10011101_01111101_11011110_11111111_11111111_11111111_11111111_00111111_01100011_11111001_11111111_11111111_11111111_11010010_01111100_10010111_11111111_11111111_11111111_11111111_00010101_01111001_11101100_11111111_11111111_10000011_11111111_11111111;
assign in[468] = 496'b11100111_10001011_11001010_11111111_11111111_11011000_01011110_01011011_01111001_10011001_11111111_11111111_01000011_00000010_00011110_01000001_01001111_11111111_11111111_01110000_01000111_01010101_11010000_01110100_11110100_11111111_01011101_00110111_11100100_11100011_01111101_11010111_11111111_11111111_11111111_11111111_11000100_01101100_11110000_11111111_11111111_11111111_11111011_01010001_10000110_11111111_11111111_11111111_11110111_00110100_01100100_11111001_11111111_11111111_11101011_01001111_01010100_11011111_11111111_01011111_11011111_11111111;
assign in[469] = 496'b11011001_01100000_01111101_01110111_11101000_11111111_00110110_01100101_00101011_01111010_11100101_11111111_11100101_01110111_10100000_00001011_01100000_11111111_11111111_10101101_01111101_11100111_00110100_00110110_11111111_11111111_00100011_00110111_11111010_01110000_00000110_11111111_11101001_01110111_10110010_11101000_01111101_10011001_11111111_11100110_01111010_10010101_10111110_01111101_10101000_11111111_11111111_00101110_01110111_00010001_01111101_01010110_11111111_11111111_11010110_01101000_01111110_01111010_11001000_11010010_10000010_10110101;
assign in[470] = 496'b01000010_00000100_11111111_11111111_11111111_11111111_00000011_00111001_11111111_11111111_11111111_11111111_11111111_10001101_01100000_11111111_11011010_11101100_11000111_00011010_01001010_01111110_00111101_01111011_00001010_11111111_11010000_00100110_01011110_11001011_11101000_11111111_11111111_11111111_00010000_00110111_11111111_11111111_11111111_11111111_11111111_00101101_00010000_11111111_11111111_11100111_11111111_11110010_01110010_10000101_10000100_00101111_01101010_11111111_11111000_01010011_01100111_00011111_10100101_11111111_11111111_11111111;
assign in[471] = 496'b11111111_11100000_01111111_11100000_11111111_11111111_11111111_00011111_01111111_01010000_11100000_11111111_11111111_00010000_01101111_00100000_01101111_01010000_11111111_10100000_01111111_10100000_11111111_11010000_01101111_11111111_01100000_01010000_11111111_11111111_11111111_01101111_10010000_01101111_11010001_11111111_11111111_11100000_01101111_01101111_10010000_11111111_11111111_11111111_10110000_01101111_00101111_11111111_11111111_11111111_11111111_00100000_00010000_11110000_11111111_11111111_11111111_11100000_01100000_11111111_11111111_11111111;
assign in[472] = 496'b11111111_11111111_01000000_11010010_11111111_11111111_11111111_10101001_00011001_11111111_11111111_11111111_11111111_11111110_01001100_11000010_11111100_11111111_11111111_11111111_10110000_01111100_01011001_01011111_10111100_11111111_11111100_01010001_10001110_11110010_11100100_00100011_11111111_10100001_01001001_11111111_11111111_10011000_10101010_11111111_00010110_00111111_11111111_11110100_00110100_11111111_11111111_11100110_01001001_11110010_00111101_10100110_11111111_11111111_11111111_00010001_01110001_10001001_11111101_11111111_11111111_11111111;
assign in[473] = 496'b11111111_10010100_01000010_11111111_11111111_11111111_11111111_10011011_00111011_11111111_11111111_11111111_11111111_11111011_01100011_10001110_11111111_11111111_11111111_11100010_00011111_01111011_01000010_00111110_11010111_11111111_11101101_01000101_01110001_00011101_11001110_11111110_11111111_11111111_01011001_00100111_11111111_11111111_11111111_11111111_11111111_01011010_10001010_11111111_11111111_11111111_11111111_11111110_01100001_10000111_10101110_10010011_00101000_11111111_11111111_00010110_01100110_00111010_00000000_11111111_11111111_11111111;
assign in[474] = 496'b10110100_01101001_01011101_00011110_11001000_11101100_01110010_10110001_11010000_10011001_01011110_11111111_11111011_01101000_10101111_11111111_11111111_10011101_11111111_11111111_00000110_00101100_11001011_00110000_01010000_11111111_11111111_11001011_01111000_01100110_11000000_11111111_11111111_11110011_00011000_01100110_00001010_11111111_11111111_11111111_00110011_00110100_11010110_01011000_11111100_11111111_10111110_01100001_11110111_11111111_00111000_10011100_11111111_10011000_01011001_11111111_10110110_00010101_10111100_01110001_00011001_10011110;
assign in[475] = 496'b11111111_11100111_01100010_11100010_11111111_11111111_11111111_00011110_10011010_11111111_11111111_11111111_11111111_11011111_01010111_11111101_11111111_11111111_11111111_11111111_00100000_01000111_00110000_00110010_11110001_11111111_11111000_01101110_00011111_11001100_00111010_10110100_11111111_00010001_00000100_11111111_11111111_01100000_11010000_11001110_01011101_11110011_11111111_10011110_00100110_11111111_11101011_10101001_11011101_10010100_01000110_11110001_11111111_11111111_10111010_01010000_01010100_11100110_11111111_11111111_11111111_11111111;
assign in[476] = 496'b11111111_11111111_11111111_11011101_10001110_11111111_11111001_10101110_00110111_01110101_01010100_10111100_00010001_01100101_01111100_01000000_11000111_11111111_00110111_00000001_01110111_00011010_11111100_11111111_11111111_11111111_10101011_01011100_11111001_11111111_11111111_11111111_11111111_00011010_00001111_11111111_11111111_11111111_11111111_11111111_00011010_00001000_11111111_11111111_11111111_11111111_11111111_10100000_01111001_00001000_10111010_10111011_10011110_11111111_11111111_10111100_00010001_01010000_01010011_11111111_11111111_11111111;
assign in[477] = 496'b11111000_01100000_11101100_11111111_11111111_11111111_10110000_00110011_11111111_11111111_11111111_11111111_11111111_00110000_10011011_11111111_11111111_11111111_11111111_11101111_01100111_11110110_10111111_00010101_10101110_11111111_10110101_00010000_10001101_01000011_10111011_01010101_11111111_00110111_00001110_01001010_11110110_11111011_01101100_11111111_01101001_01100010_11100111_11111111_10010011_01000101_11111111_00110101_10011001_11101011_10010000_01010000_11110001_11111111_11111111_10111010_01110001_00100111_11101011_11111111_11111111_11111111;
assign in[478] = 496'b00101011_01111011_01000001_11111111_11111111_11100001_01110101_01110111_10100001_11111111_11111111_11111111_00010000_00111010_10110011_11111110_11111111_11111111_11110010_01111000_10110011_11111111_11111111_11111111_11111111_10111011_01100110_11110001_11111111_11111111_11111111_11111111_11000101_01101010_11101011_11111111_11111111_11111111_11111111_11110100_01110001_00100000_11111010_11111111_11111111_11111111_11111111_11010101_01011101_00000111_10101001_00001101_01001000_11111111_11111111_11011011_01011010_01111101_01000110_11111111_11111111_11111111;
assign in[479] = 496'b11111111_11010000_00011111_01011110_01111100_11011000_00010101_01011010_10110101_11100100_11100100_00000110_01010100_10010100_11111111_11111111_11111111_11101011_00101011_11111000_11111111_11111111_11111111_11111111_10100000_11111001_11111111_11111111_11111111_11111111_11011001_01011110_10011000_11111111_11111111_11111111_11111111_00011000_00110011_01100001_11111101_11111111_11111111_10100010_01011101_11100101_00111001_00000010_11111010_10100010_01011100_11001000_11111111_11010001_01110101_01001001_01011100_10110101_11111111_00101111_11001100_11111111;
assign in[480] = 496'b01111000_00110101_00000111_01001010_10011011_01011100_11001100_11111111_11111111_11111111_11111111_01110000_11011111_11111111_11111111_11111111_11111111_11111111_01100000_00110100_11011000_11101110_11111111_11111111_11111111_11100100_00110101_01111101_01101011_10001001_11111111_11111111_11111111_11111111_10110001_01111101_01001100_11111111_11111111_11111111_11100010_01101010_01001010_11001111_11111111_11111111_11111111_10100001_01111100_01011001_00000110_10010100_10010101_11111111_11111001_10011001_00100110_01111000_01111110_11111111_11111111_11111111;
assign in[481] = 496'b01011111_10110010_11111111_11111111_11111111_11111011_01100100_10110010_11111111_11111111_11111111_11111111_11100010_01111101_11101010_11111111_11111111_11111111_11111111_11010011_01111110_11101110_11111111_11111111_11111111_11111111_10100110_01001010_11111100_11111111_11111111_11111111_11111111_00010100_00011111_11000001_11111111_11111111_10000010_11111001_01011111_00101101_00111011_00110010_11101010_11001101_11101110_01010011_11111111_11111100_10100010_01001101_00100000_11111100_11010101_11111111_11111111_11111111_11101001_11111111_11111111_11111111;
assign in[482] = 496'b11111111_10101011_01001101_00100001_00101100_11111111_11111010_01010110_11011111_11010100_00110010_11111111_11111111_10110101_00001011_11100001_01000011_11000110_11111111_11111111_10011111_00111011_01001100_11000111_11111111_11111111_11111111_10000001_01001110_11111000_11111111_11111111_11111111_10001110_01101101_00110000_11111111_11111111_11111111_10111011_01011010_11010111_01001011_11111110_11111111_11111111_00010110_00100110_11101000_00001010_11101010_11111111_11111111_11101000_10000111_01001101_01001010_11011000_11111111_10110110_10001111_11111111;
assign in[483] = 496'b11111111_11111111_00100000_10110110_11111111_11111111_11111111_10010011_10011101_11111111_11111111_11111111_11111111_11011011_00110010_11111110_11111111_11111111_11111111_11111110_00101101_11011111_11111111_11111111_11111111_11111111_10101010_10001011_11111111_11111111_11111111_11111111_11111111_00111010_11110100_11111111_11111111_11111111_11111111_11101010_00010110_11111111_11111111_11111111_11111110_10101111_11101010_00110010_11101100_11001110_10001001_00001100_10110100_11111111_10110110_10000110_10010000_11011111_11111111_11111111_11111111_11111111;
assign in[484] = 496'b11111111_11111111_11001110_01100001_00001001_11111111_11111111_11100000_01101001_00101011_11111011_11111111_11111111_11101101_01001011_00110111_11111100_11111111_11111111_11111010_00101110_01001011_11111011_11111111_11111111_11111111_10011010_01101110_11011110_11111111_11111111_11111111_11101110_01101111_10101101_11111111_11111111_11111111_11111111_10100010_01100000_11111110_11111111_11111111_11111111_11111111_11001101_01110010_10110111_11010111_10111110_00011100_00000111_11111111_00010101_01101111_01111110_01100101_00100110_11111111_11111111_11111111;
assign in[485] = 496'b11111111_11111111_10101111_01101001_11001101_11111111_11111111_11001110_01110011_10111001_11111111_11111111_11111111_11111111_01001011_00000100_11111111_11111111_11111111_11111111_10100101_01011111_11101100_11111111_11111111_11111111_11110110_01001011_10111001_11111111_11111111_11111111_11111111_10011011_01010101_11110110_11111111_11111111_11111111_11111111_00110111_10111001_11111111_11111111_10101111_11111111_11110110_01011111_11010111_11001101_00001110_01001011_11110110_11111111_00101100_01111101_01001011_10010000_11101100_11111111_11111111_11111111;
assign in[486] = 496'b11111000_01000011_01101011_00110011_11111111_11111111_00001001_00001010_11111100_00111111_11111110_11111111_11111111_01001001_11011101_11101001_01001111_11111111_11111111_11111111_10000101_10011011_00110011_10010101_11111111_11111111_11111111_10110011_01111000_00011000_11111110_11111111_11111111_11001111_01010110_01110010_11001100_11111111_11111111_11111111_00110011_11000011_10110010_00111001_11111111_11111111_11111111_11111010_11111101_11111111_01000110_11001010_11111111_11111111_11111000_10001101_11111111_00100100_11001001_00110010_01010100_01001000;
assign in[487] = 496'b11000001_01000100_01011011_11000001_10110100_11101011_01010111_00010001_00000111_01010100_00100010_11111111_10100010_01000000_11111110_11111111_11111111_11111111_11111111_00001000_00010000_11111111_11111111_11111111_11111111_11111111_10110110_01110100_10010111_11101001_11111111_11111111_11111111_11111100_10100001_01100101_01000101_11111111_11111111_11111111_11111111_11110010_01001010_10000100_11111111_11111111_11111111_11011010_01011010_00110011_11111111_11111111_11111111_11111111_00000111_01111101_11000101_10101110_00110110_00001111_01100001_01101010;
assign in[488] = 496'b11111111_11111111_00000000_00100110_11111111_11111111_11111111_11111111_01010011_10100010_11111111_11111111_11111111_11111111_10111101_01110110_11011100_11111111_11111111_11111111_11111110_00100101_01011100_00101010_11111111_00010111_00111001_01101001_01111110_00100110_11100001_11111111_11011010_11011010_00101110_00100110_11111111_11111111_11111111_11111111_11100111_01111010_00000100_11001001_11111100_11111111_11111010_01001100_01100111_01000001_01110001_00111010_11100111_11100001_00101010_11111100_11111111_11101001_00001001_11111111_11111111_11111111;
assign in[489] = 496'b11111111_11111111_11011100_00001001_01110011_11111111_11111111_10001100_01110101_01111110_01011101_11111111_11111111_10101011_01110111_00101000_10111111_11111011_11111111_11111111_00010111_01011001_11101010_11111111_11111111_11111111_11111111_00000011_01111110_01000100_11111111_11111111_11111111_11111111_11101000_01100000_01100010_11111111_11111111_11111111_11111111_10101100_01111011_00100110_11111111_11111111_11111111_11100101_01110111_01010001_11000111_11111111_11111111_11111111_11001111_01111110_01110001_01010100_11111111_00011111_01010101_10001010;
assign in[490] = 496'b11111111_11111111_11101111_01111100_01111011_11111111_11111111_11111111_10001110_01111101_01001001_11111111_11111111_11111111_11000011_01010100_01100011_10111111_11111111_11111111_11100010_01001100_01111011_00100010_11111111_11111111_11110110_00010010_01111101_01011011_11001111_11111111_11111111_00001110_01111011_01101101_11000001_11111111_11111111_10111111_01100010_01111100_10000111_11111111_11111111_11111111_01001001_01111011_00010011_11111111_11111111_11111111_11111111_01001001_01101100_10110001_11111111_11111111_11111111_11111111_11111111_11111111;
assign in[491] = 496'b11111111_11111111_10000010_01111100_10100000_11111111_11111111_11110100_01011001_01111101_10001100_11111111_11111111_11111111_00110111_01111011_01111100_11111111_11111111_11111111_11110101_01100000_01111011_10101011_11111111_11111111_11111111_00110000_01111101_01110100_11011100_11111111_11111111_11100010_01110001_01111100_10100011_11111111_11111111_11111111_00101000_01111100_01110001_11011101_11111111_11111111_10101101_01111011_01111011_10011011_11111111_11111111_11111111_00100001_01111011_00000100_11111110_11111111_11111111_11111110_11111111_11111111;
assign in[492] = 496'b11111111_11100000_10100000_00000000_11100000_11111111_00010000_01111111_01111111_01111111_01101111_11110000_01010000_01111111_01100000_11110000_11110000_00101111_00011111_01111111_01101111_10110000_11111111_11111111_00000000_01111111_01101111_11000000_11111111_11111111_10110000_01111111_00010000_11010001_11111111_11111111_11010001_01111111_01010000_11111111_11111111_11111111_11010000_01101111_01111111_11110000_11111111_11111111_11000000_01101111_01101111_11010001_11111111_11111111_11000000_01101111_01010000_11010001_11111111_01111111_11010001_11111111;
assign in[493] = 496'b11111111_11111111_11111111_11111111_11111111_00010110_11010110_11111111_11111111_11100001_00000101_11001011_01111101_11001110_11101110_00010100_01110011_01001100_11100110_01111101_10011010_01100110_01110011_10011100_10101101_11110010_01101110_01111101_01111101_01011011_01111001_01111101_10100010_01110111_00101110_00011101_00011101_00010000_10110000_01101110_10001100_11111111_11111111_11111111_11111111_11111111_01110000_11110001_11111101_11111010_11111111_11111111_11111111_01111001_00011110_01001011_00100100_11111111_11111111_01011010_11000110_11111111;
assign in[494] = 496'b10000011_01010001_11110001_11111111_11111111_11111110_01000001_11011000_11111111_11111111_11111111_11111111_10101110_00011000_11111111_11111111_11111111_11111111_11111111_01000011_11001010_11111111_11111111_11111111_11111111_11110100_01010001_11111000_11111111_11111111_11111111_11111111_11011011_00110011_11111111_11111111_11111111_11111111_11111111_11110010_01100011_11001011_11111111_11111111_11111111_11110111_11111111_10110110_01000111_00111011_10000011_10011010_01010111_11111111_11111111_11111111_11011001_10000011_10000001_11111111_11111111_11111111;
assign in[495] = 496'b11111111_11111111_11111111_11111111_11111111_00011110_01101100_01111100_01001011_10100001_11111111_01101010_00010101_10111111_10111111_00010101_01111001_00001110_10110011_11111111_11111111_11111111_11101111_01100110_01110110_11110110_11111111_11111111_10111100_01010011_00001111_01100111_01011100_00011011_01000001_01111010_00001011_11101101_01101011_00011110_00110101_00001010_11010101_11111111_11001001_01111010_11111111_11111111_11111111_11111111_11111111_01001101_00010111_11111111_11111111_11111111_11111111_10111110_01101010_11111111_11110000_01001101;
assign in[496] = 496'b11110010_00101101_01111101_01111101_01111001_11111111_10110001_01111011_00001111_11010101_00101101_11111111_11111111_11001101_01110001_10111001_11111000_01010101_11111111_11111111_11111111_00011001_01011110_00111101_01110000_11111111_11111111_11111100_10010111_01111110_01111110_10011010_11111010_10011110_01101011_01111101_01110101_01111101_10101010_00111110_01111101_01001100_10101010_11011010_01101100_10001110_01011011_01100101_00101111_11010100_00100111_01111101_10110101_11011001_10001001_01111110_01111101_01111000_00011001_11000000_10000100_11000100;
assign in[497] = 496'b11011010_00100010_01011111_01101111_00010110_10010000_01010011_10011111_11110010_11011111_00110101_00000100_00100100_11110001_11111111_11111111_11111111_11000000_00110001_11111100_11111111_11111111_11111111_11111111_11011001_11000000_11111111_11111111_11111111_11111111_11111111_10011011_11111100_11111111_11111111_11111111_11111111_11111111_00110001_11111100_11111111_11111111_11111111_11111111_10111101_01000001_11000000_11111111_11111111_11111111_11111010_01011111_11000000_01010000_10101101_00000101_10001101_00111000_10001011_11010011_01001000_10011100;
assign in[498] = 496'b11111111_11111111_11111111_11111111_11111111_11110110_10100011_01001110_01011110_00000110_11111111_11110011_00111001_00000000_11100110_11101111_01000101_11011011_00010101_11011010_11111111_10000011_10010101_00011010_10111110_00111001_10010111_00010101_10011001_11110111_00101110_11110011_10011100_10011110_11111100_11111111_11010010_00101000_11111111_11111111_11111111_11111111_11111111_00011100_10111111_11111111_11111111_11111111_11111111_11110101_00110000_11111111_11111111_11111111_11111111_11111111_10011110_00010001_11111111_11111111_00111111_11100111;
assign in[499] = 496'b11111111_11111111_11111111_11111111_11111111_11111110_11111000_11111111_11111111_11111111_11000101_01001000_01110010_00111101_11011101_00000100_01101010_01111101_10011001_10001010_01111100_01111101_01111100_01011011_10010000_11110110_00111101_01111101_01100011_01111101_01111101_01111110_00111011_01111010_10001110_11111111_11010100_10010101_11000100_01111000_10010011_10110111_00000010_11111111_11111111_11111111_01111101_01110110_01111101_01110110_11110011_11111111_11111111_00011001_00100001_00000100_11110001_11111111_11111111_11111111_11111111_11111111;
assign in[500] = 496'b10011101_01000100_01110111_00111011_10101101_01000110_01010010_10100010_11000101_10010110_01100110_00010001_00011000_11110001_11111111_11111111_11111111_00110111_01101001_11110010_11111111_11111111_11111111_11111111_00110111_01000100_11111111_11111111_11111111_11111111_11100011_01101010_01101010_11111111_11111111_11111111_11111111_00001000_01100101_00101101_11000111_11111111_11111111_11011101_01110011_10110011_11011001_00111101_11111101_11100001_01010000_00011001_11111111_11111111_00111001_01001000_01100010_00010110_11111111_01001111_10110011_11111111;
assign in[501] = 496'b11111111_11111100_10000011_01101001_01111101_11111111_11111111_10101110_01110110_00000110_00000011_11111111_11111111_11111111_00000111_00111101_11011011_00101100_11111111_11111111_11111111_00100100_01110001_01110101_01101111_11111111_11010110_01000111_01111101_01111100_10000001_11111000_10001100_01101101_01011000_01000110_01011010_11111111_11111111_01111101_00010111_11111000_00101000_00100111_11111111_11111111_01011011_11111001_11101011_01101010_10101001_11111111_11111111_01010111_00010101_01110000_01000101_11111110_11111111_00010011_11101001_11111111;
assign in[502] = 496'b11111111_00100110_10100110_11110010_00111001_11111111_11111111_11001010_00111011_00101101_10001101_11111111_11111111_11111101_10010001_01111110_10010111_11111111_11111111_10111001_01010000_00001010_00011100_10001110_11111111_11001010_01100111_11010001_11111111_11011010_00111111_11111111_00101111_10110100_11111111_11111111_11111111_01010000_11111111_01010000_11111111_11111111_11111111_11010111_01000100_11111111_00101100_10101000_11111111_11111111_10001000_10110000_11111111_11101011_00011111_01000010_00001110_00101001_11111110_11110001_10011111_11111011;
assign in[503] = 496'b11111111_11010010_01111101_00111100_11111111_11111111_11111111_01000000_01111110_10101110_11111111_11111111_11111111_10100100_01111100_00100000_11111111_11111111_11111111_11101111_01101101_01100101_11110010_11111111_11111111_11111111_00100101_01111101_10010111_11111111_11111111_11111111_11110111_01111000_01101001_11110100_11111111_11111111_11111111_11111000_01110101_00100111_11111111_11111111_11111111_11111111_11111111_10101000_01101011_10000111_10100001_11001111_11111111_11111111_11111111_11100100_10100100_00111011_01001011_11111111_11111111_11111111;
assign in[504] = 496'b01011011_10100100_11111111_11111111_11111111_11111111_01001001_10100011_11111111_11111111_11111111_11111111_11111111_01110110_11000110_11111111_11111111_11111111_11111111_11111111_01000100_11000011_11110001_00101101_01000000_11111111_11111111_01111101_11011001_00111110_01111001_00111111_11111111_11111111_01111000_00011101_00111001_01011000_00000000_11111111_11111111_01010100_01110010_10010000_01110010_11101100_11111111_11111111_01000011_01110101_01100110_10110011_11111111_11111111_11111111_00110111_01001111_11001111_11111111_11111111_11111111_11111111;
assign in[505] = 496'b11111111_11111111_11111111_11111111_11111111_01101111_11111111_11111111_11111111_11111111_11111111_00010000_01111111_11110000_11111111_10110000_10100000_11110000_00000000_01111111_00100000_01100000_01111111_01111111_01111111_00000000_01111111_01111111_00101111_11010000_11111111_01010000_00100000_01111111_00000000_11111111_11111111_11111111_00100000_01000000_01010000_10010001_11111111_11111111_11010001_01101111_11010000_11100000_01101111_00100000_00010000_01101111_01100000_11111111_11111111_10110000_01101111_01101111_00010000_11111111_11111111_11111111;
assign in[506] = 496'b00111000_10011011_11000101_01001001_11111111_00111011_11100110_11111111_11101100_00110010_11111111_11111111_00110100_11111110_11111111_00000011_10110100_11111111_11111111_00001001_10111101_11011011_00010001_11111111_11111111_11111111_11110001_01000100_00111101_11111000_11111111_11111111_11111111_11111111_00101011_01000011_11011000_11111111_11111111_11111111_10000100_10110000_11100101_01000110_11010000_11111111_11101110_10110011_11101111_11111111_11100110_00100101_10101001_11111111_11111111_00110110_10100001_10110011_10111111_11010010_10011101_10011101;
assign in[507] = 496'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111110_11010000_10011111_10011010_11111111_11111111_11011000_00111101_10001010_10110001_11000001_11111111_11111111_11101010_00010001_11000100_11111111_11111111_11111111_11111111_11111111_11111011_10101011_00011100_11000101_11111111_11111111_11111111_11100111_10000001_00101011_10101001_00010000_00111010_01001101_00111010_10010010_11010001_11111111_11000110_11101111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111;
assign in[508] = 496'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_11100100_10001111_00101011_00010101_11111111_11111111_10011101_01110001_01111111_01111111_01111111_11111111_10111001_01111111_01100011_10001111_10111001_10101011_11111111_10010110_01111111_10001000_10111010_11100100_11111111_11111111_11111111_00111000_01111111_01110001_10111001_11111111_11111111_10101011_01100011_00100011_11100100_11111111_11111111_01011100_01011100_00000000_11110010_11111111_11111111_11111111_10111001_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111;
assign in[509] = 496'b11111111_10111100_01110010_00110010_11111111_11111111_11111111_10011010_01111011_10011000_11111111_11111111_11111111_11101100_01100101_01000011_11111111_11111111_11111111_11111111_00011110_01111101_10100010_11100001_11100001_10100011_01101000_01111100_01111110_01111101_01111101_01111101_11001001_01111011_10010101_11100000_11100000_01001111_01100101_00010011_00110000_11111110_11111111_10011110_01110010_10110111_01101011_11010100_11111111_10101010_01110110_10001001_11111111_00001011_11111111_11111111_00101111_10000011_11111110_11111111_11111100_11111111;
assign in[510] = 496'b01001000_11111111_11111111_11111111_11111111_10110110_01111100_11110110_11111111_11111111_11111111_10010010_01011111_01111111_11110010_11111111_11111101_00011111_10011010_01010111_01111110_01101111_01011000_01101100_01111110_11111111_11000101_01111110_10110111_10100110_10110110_01000111_11111111_11000101_01111110_11110101_11111111_11111111_01000011_11111111_11000101_01111110_11110101_11111111_11111111_01000011_11111111_11000101_01111110_11110101_11111111_11111111_00111000_11111111_11101011_01111110_10110100_11111111_11111111_00010010_10010110_11111111;
assign in[511] = 496'b11111111_11111111_11111111_11111111_11111111_11111110_10111011_00001010_00101011_01111000_01101010_11111111_10100011_01111100_01111101_01100010_00011011_01001110_00001110_01111010_01111101_01010111_11110001_11111110_00110110_01111101_01111100_01010000_11010111_11111111_00000101_01111100_01111110_00000101_11110000_11111111_10011111_01111100_00011010_11100110_11111111_11111111_10101111_01110010_00111001_11111111_11111111_11111111_10101010_01111001_00101011_11110000_11111111_11111111_10101100_01111011_01010100_11011010_11111111_01000101_11111100_11111111;
assign in[512] = 496'b01111011_01111011_01111100_01100100_10010001_01001110_10111110_11110110_11110110_11010101_00101001_01111011_10010101_11111111_11111111_11111111_11111111_11110111_01001111_00110111_11110011_11111111_11111111_11001111_10000110_11101011_00110010_01011111_00111010_01100000_01110100_01100001_11111111_11111111_00100110_01111011_00101111_00000011_11111110_11111111_10011011_01111000_10001110_11111111_11111111_11111111_11111111_00010000_01010001_10010110_11101100_11010110_10000100_11111111_10111011_01101110_01111011_01111100_01111011_11101001_11001001_10000001;
assign in[513] = 496'b11111111_10111010_01111101_11110010_11111111_11111111_11111111_10101101_01101011_11111000_11111111_11111111_11111111_11111111_00011110_00101000_11111111_11111111_11111111_11111111_11110111_01101101_10001010_11111111_11111111_11111111_11111111_00001000_01010100_11101010_11111111_11111111_11111111_11000010_01111001_10101100_11111111_11111111_11111111_11111111_00110001_01101011_10101001_10010011_10000011_00000011_11111111_01001011_01111110_01001001_00111001_01000011_00100011_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111;
assign in[514] = 496'b11111111_11100011_10011000_10110000_11111011_10010110_00111100_01110100_01110000_01101101_00101100_11111111_00010001_01111110_00111110_11101001_10010011_01110100_11000011_01111101_01111101_10101010_11111111_01000110_01100111_00111011_01111101_01011100_11111100_10101001_01111110_10010001_00010110_01110101_10110100_11101000_01100001_01010111_11111011_11111100_11110001_11111111_00010011_01110111_11000111_11111111_11111111_11111111_11101000_01110111_00101000_11111111_11111111_11111111_11111110_00111001_01111101_11011010_11111111_01111101_00000111_11111111;
assign in[515] = 496'b01111110_01111010_01101011_01101001_11011000_11001010_01101100_11011110_11110111_01011100_00111000_11111111_11111000_01110001_10111001_11111101_01100010_01010101_11111111_11111111_10010001_01011100_00011010_01111110_00010000_11111111_11111111_11110111_01101010_01111110_01010001_11110010_11111111_11101110_00111010_01111110_01111100_11010000_11111111_11001101_01011110_01110011_00100101_01111110_11001000_11111111_01111010_01011001_00111001_11010010_01111010_10001111_11111111_00101011_11101010_00001111_01111000_01111101_10110011_11111101_10101010_10111010;
assign in[516] = 496'b11111111_11111111_11010001_01111111_01000000_11111111_11111111_11111111_00100000_01111111_10110000_11111111_11111111_11111111_11000000_01111111_01010000_11111111_11111111_11111111_11111111_01000000_01111111_11000000_11111111_11111111_11111111_11000000_01111111_01000000_11111111_11111111_11111111_11111111_01000000_01111111_11010001_11111111_11111111_11111111_11010001_01111111_00100000_11111111_11111111_11111111_11110000_01010000_01111111_11100000_11111111_11111111_11111111_00000000_01111111_00011111_11111111_11111111_11111111_11111111_11111111_11111111;
assign in[517] = 496'b11111111_11111111_11000111_00010011_10010010_11111111_11011111_00101101_01111001_01111010_01100010_11111111_11010010_01101001_01100010_10010011_11100010_11111111_11111111_00101010_01011011_11110001_11111110_11111010_11111111_11111111_10110011_01110010_00101001_01011100_01011010_11111100_11111111_11001111_01100100_01100100_00101001_10010001_11111111_11000101_01101100_00110101_11100110_11111111_11111111_11111111_01000011_00111011_11111101_11111111_11110000_11111110_11111111_01010011_00101111_00010011_01001111_01110110_11000010_00111101_00010101_10101100;
assign in[518] = 496'b01110101_11100100_11111111_11111111_11111111_00010000_00111111_11111111_11111111_11111111_11111111_11111111_00010001_00010001_11111111_11111111_11111111_11111111_11111111_00010000_00101010_11111111_11111111_11111111_11111111_11111111_00010001_01101011_11101110_11111111_11111111_11111111_11111111_10100011_01111100_10001111_11111011_11111111_11111111_11111111_11111111_00010000_01111101_00101100_11001010_11101001_11111111_11111111_11111110_00100011_01110010_01111101_01110010_11111111_11111111_11111111_11111111_11101001_11001010_11111111_11111111_11111111;
assign in[519] = 496'b11111111_11111111_00011011_01101100_11101110_11111111_11111111_10100100_01111101_10100110_11111111_11111111_11111111_10110100_01111000_00111010_11111000_11111111_11111111_00011100_01101110_01111101_01011000_00101110_00100001_11111111_01011000_01111011_10010001_10101110_10010100_01111000_11100101_01111000_00010111_11111111_11111111_10010100_01110100_10011110_01111011_11001010_11111111_10101111_01110010_10100011_00010011_01000110_11111111_11111111_00100110_00011000_11111111_10001111_00111001_11111111_11111111_11111101_11111100_11111111_11111111_11111111;
assign in[520] = 496'b01011101_10101101_11111111_11111111_11111111_10100001_01110100_11101111_11111111_11111101_10011100_11111111_10000010_01010011_11111111_11011010_01000010_01111100_11111111_11001101_01111000_00101111_01110010_01111101_01111101_11111111_11111111_00110001_01110101_00111110_00011001_10110010_11111111_10000010_01111101_10100000_11111111_11111111_11111111_11010111_01110111_00011110_11111101_11111111_11111111_11111111_00001000_01110101_11101100_11111111_11111111_11111111_11111111_00010100_01001110_10001010_01010001_01110010_11110011_01100111_00001010_11101111;
assign in[521] = 496'b11111111_11111111_11111111_11111111_11111111_11111111_11110101_10111111_10110110_10000111_10101010_11111111_11000011_01101000_01101001_01010010_01010010_01000110_11110110_01101110_00010011_11110100_11111111_11111111_11111111_11111111_00110011_10011001_11001000_11000110_11111111_11111111_11111111_10010001_01111101_01111101_01111001_11110010_11111111_11100100_01101101_01100000_10010101_10011111_11101011_11111111_10101100_01111101_00111011_01000000_01111101_10001010_11111111_11111111_10001100_00110001_00110001_10010000_11111001_11111111_11111111_11111111;
assign in[522] = 496'b11111111_11111111_01011010_00001111_11111111_11111111_11111111_11111111_01101110_00011111_11111111_11111111_11111111_11111111_11010101_01111010_10011111_11111111_11111111_11111111_11111111_10010010_01101010_11110010_11111111_11111111_11111111_11111001_01100100_00100111_11111111_11111111_11111111_11111111_11110011_01111101_10011000_11111111_11111111_11111111_11111111_10110001_01111010_11101011_11111111_11111111_11111111_11111111_00011010_01000110_11111111_11111111_11111111_11111111_11101000_01100111_00001111_11111111_11111111_01000011_11110111_11111111;
assign in[523] = 496'b11111111_11100000_11010011_11011111_11111111_11100100_01001001_01110111_01110010_01110011_01000010_11111111_00000100_00110011_11101111_11111111_11111110_10011111_11111111_11100000_01001101_10010001_11100110_11111111_11010010_11111111_11111111_11100000_00001000_01011001_01010101_10001001_11111111_11111111_11111111_11111101_10000100_01111110_01001011_11111111_11111111_11111101_00000100_01101111_10100000_11111000_01000010_01000010_01010001_01111110_11001011_11111111_11111111_10100011_10100011_10100011_11010100_11111111_11111111_11111111_11111111_11111111;
assign in[524] = 496'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_11000010_10001001_00101001_00101001_11111111_10000100_01110000_01110001_00110101_00010000_00000011_11101000_01111010_10100101_11100100_11110100_11111111_11111111_11101110_01110100_00101011_01101010_01001000_11111111_11111111_10111011_01110100_01101010_00101100_10110101_11111111_11111111_01110000_00101100_11110100_11111111_11110001_11001011_11111111_00100101_00111001_10010000_10001111_01010001_01101011_11111111_11100111_00100011_01100001_01100001_00101111_11001110_11111111_11111111_11111111;
assign in[525] = 496'b11101011_01101111_01100111_00111110_01110111_11111111_11000000_01001100_11111011_10101000_01111101_11111111_11111111_10101100_00110100_11001000_01110100_00001101_11111111_11111111_11001001_01110110_01110010_00111110_11111110_11111111_11111111_10001110_01111110_00111111_11111000_11111111_11111111_00000101_01111011_01101100_00110111_11111111_11111111_10010010_01111101_00001011_10110011_01010100_11111111_11111111_01111101_01001100_11110111_00001000_01110010_11111111_11111111_01101000_01111100_01110100_01111101_00101101_11111111_10000010_11000001_11111110;
assign in[526] = 496'b11111111_11111111_11111111_11000111_01011001_11111111_11111111_11111111_10000001_01111011_01111100_11111111_11111111_11111111_11110001_01010100_01111100_00111010_11111111_11111111_11111111_10001111_01111011_01001110_11101000_11111111_11111111_10110100_01111110_01010011_11110111_11111111_11111111_10001110_01111100_01100001_11011010_11111111_11111111_11000100_01110010_01101110_11010100_11111111_11111111_11111111_01010111_01111010_10100101_11111111_11111111_11111111_11111111_01111100_10001010_11111111_11111111_11111111_11111111_11111111_11111111_11111111;
assign in[527] = 496'b11111111_11111111_11111111_11111111_11111111_11000100_01000010_01100101_01000111_11100111_11111111_11100101_00110100_10110110_00000111_00101001_00100111_11111111_11110001_01000000_01100000_10111000_11111000_00111110_11111110_11111111_11111111_11111111_11111111_11111111_01010100_11100111_11111111_11111111_11111111_11111111_11111111_01010011_11110110_11111111_11111111_11111111_11111111_10011010_00000101_11111111_11111111_11111111_11111111_11111110_01010000_11101011_11111111_11111111_11111111_11111111_00000101_10011001_11111111_10111010_00110111_11111001;
assign in[528] = 496'b11111111_11110101_10010001_10000110_11010101_11111111_11111111_00010101_01111111_01111110_01111111_11111111_11111111_11111111_01011100_01111110_10111111_10001010_11111111_11111111_11111111_01000111_01111110_01001110_10101101_11111111_11111111_11110110_01000011_01111110_01111000_10010110_11111111_11100100_10001010_01111110_01100101_10001101_11111111_10001010_01110101_01111110_00100111_11111000_11111111_11111111_01111111_01001100_00000101_11011111_11111111_11111111_11111111_00001100_11111100_11111111_11111111_11111111_11111111_11111111_11111111_11111111;
assign in[529] = 496'b00101100_11111111_11111111_11111111_11111111_00011111_10011111_11111111_11111111_11111111_11111111_11111111_01011110_11000101_11111111_11111111_11111111_11111111_00010110_01111100_00110010_00110001_00001100_10000111_10111000_00010111_00110011_11001011_11010001_10010010_00011111_01011110_00101111_10110101_11111111_11111111_11111111_11111111_11001000_01111010_11111111_11111111_11111111_11111111_11100001_01100001_00101100_11111111_11111111_11111111_11111111_10101100_01100100_11011110_11111111_11111111_11111111_11111111_10010011_11111111_11111111_11111111;
assign in[530] = 496'b11111111_10011111_01111011_01111011_01111011_11111111_11111101_00010010_01111011_01111011_00110011_11111111_11111111_11011010_01111100_01111011_01110110_11001010_11111111_11111111_10100110_01111100_01111011_01101001_11111111_11111111_11111111_00000111_01111101_01111100_10000111_11111111_11111111_11111111_01000010_01111100_01111011_11011001_11111111_11111111_10111111_01111000_01111100_01001011_11111010_11111111_11111111_10010110_01111011_01111100_10000001_11111111_11111111_11111111_00011111_01111011_01111100_11111001_11111111_01001000_00110010_11111111;
assign in[531] = 496'b10101100_00010011_00110110_00110110_11001010_01010001_01110100_01001100_00010101_01100100_01101100_01110100_00011010_11101010_11111111_11111111_11111111_00110110_00101011_11111111_11111111_11111111_11111111_11111111_11010111_11101101_11111111_11111111_11010010_10100110_11111111_11111111_11111111_11111111_11111111_10010110_00000111_11111111_11100010_11111111_11111111_11111111_00101100_10100100_11111111_00000011_10011101_11111111_11110011_01111110_10110101_00011001_01011001_01101100_00111011_01000000_01111101_01010101_00111111_00110011_10001111_11001010;
assign in[532] = 496'b11111001_10101100_01101010_01011010_11011100_11101010_00010001_01000101_10111000_10001101_00110001_00010110_01111000_01110111_10100011_10101100_00111011_01000100_11111010_01100110_00100000_00101111_00010000_00001101_11011001_10111011_01010110_11111101_11111111_11111111_11111111_11111111_10010101_10001011_11111111_11111111_11111111_11111111_11111111_10010101_00000010_11111111_11111111_11111111_11111111_11111111_10111010_00111101_11111101_11111111_11111111_11111111_00010000_11111101_00110110_00010000_11011011_11100001_00111011_00001010_01110100_01111011;
assign in[533] = 496'b11111111_00101011_01010101_11111011_11111111_11111111_11001101_01111010_10010110_11111111_11111111_11111111_11111111_00001110_01011010_11111010_11111111_11111111_11111111_11110011_01110001_10001111_11111111_11111111_11111111_11111111_10111001_01111011_11000111_11111111_11111111_11111111_11110110_01001010_01010000_11111111_11111111_11111111_11111111_10000100_01111101_01100110_00010010_10001011_10111101_11110110_11110110_10110000_10001001_00010100_00111110_01110110_01101001_11111111_11111111_11111111_11111111_11111111_11101001_11111111_11111111_11111111;
assign in[534] = 496'b10010010_01100110_01111110_01011001_11001101_00010101_01111110_01111110_01111110_01111110_10001101_11111111_00100101_01111110_01011101_01111110_01111100_11000100_11111111_11101101_01001011_01111111_01111110_10000011_11111111_11111111_11111111_00100000_01111110_01111110_00011101_11100101_11111111_11111111_00100110_01111110_01111110_01111110_01000011_11100010_11111010_10110011_00010111_10100011_01111110_01110101_00110000_00111001_10011000_01100110_01111110_01111110_00000111_10001110_01111110_01111110_01111110_01001100_10110000_00100100_10110011_11111111;
assign in[535] = 496'b10101010_01010101_01101010_00011000_10000110_10010111_01100111_10111001_11111001_11111111_11111111_11111111_01100000_00000101_11111111_11111111_11111111_11111111_11111111_00101001_01000111_11111111_11111111_11111111_11111111_11111111_11000010_01101101_01000010_10101110_11110110_11111111_11111111_11111111_11100111_00011111_01111101_10000101_11111111_11111111_11111111_11110110_01011101_00011000_11111111_11111111_11111111_11111111_10010101_01101011_11111110_11111101_11011100_11111111_11111111_00001001_01111101_01011110_01011010_11101110_10001100_10000001;
assign in[536] = 496'b11101110_10100101_10000010_11001100_11111111_00010100_01101011_01111101_01111100_01111001_00100100_00011100_01111101_01111101_01111110_01111101_01111110_01111101_01111101_01010011_10110110_10101001_01111100_01111101_01111100_01111101_11001111_10011001_01101111_01111100_01111101_01100011_01111110_01001110_01111101_01111110_01111101_01111110_00110100_01000010_01000010_00010111_10010010_01111100_01111101_11010101_11111111_11111111_11111111_10010110_01111101_01000011_11111111_11111111_11111111_11111111_00011110_01111100_11000010_11111111_01000001_01101100;
assign in[537] = 496'b00101011_01111101_00101010_11111111_11111111_11101011_01011011_01111110_10001001_11111111_11111111_11111111_11011001_01111011_01111101_11000011_11111111_11100001_11111111_01000110_01111101_00010100_11111110_10110010_01110001_10000111_01111100_01011111_11011101_11110100_01010010_01111100_01110000_01111100_01100000_11010000_00001001_01111101_01100011_01111110_01111101_01111101_01111110_01111101_01111110_10101010_10111111_11110010_00011000_01111101_01111100_01011010_11011001_11111111_11111111_11110010_00010011_01110101_10011011_11111111_11111111_11111111;
assign in[538] = 496'b10011111_01100011_11111111_11111111_11111111_11111111_10011111_01001001_10110010_11101110_11111111_00010110_00101000_01010101_01110101_00011011_11010111_11111111_11101111_11011100_00101001_10010100_11111111_11111111_11111111_11111111_11111111_01010101_10111111_11111111_11111111_11111111_11111111_11111110_01100100_11001011_11111111_11111111_11111111_11111111_11111011_01111101_11010110_11001111_10111010_10100011_11111111_11111101_01101100_01111100_01111100_01111101_01011100_11111111_11111111_11001000_10101111_11001010_11100010_11111111_11111111_11111111;
assign in[539] = 496'b01011110_00011110_00110101_11111010_11111111_01010001_11110000_11111111_11111111_11111111_11111111_11101000_01001111_11100011_11111111_11111111_11111111_11111111_11111111_10110111_01000000_11101110_11111111_11111111_11111111_11111111_11111111_10111111_01000010_11010010_11111111_11111111_11111111_11111111_11111111_11011100_01011011_11111000_11111111_11111111_11111111_11111111_11100100_01101001_11110011_11111111_11111111_11111111_11010010_01011101_10101110_11111111_11111111_11111111_11111111_00100101_00010010_11100100_11000110_11111011_10110111_10000001;
assign in[540] = 496'b11111111_10000010_01111100_10101101_11111111_11111111_11111111_00101100_01111100_00011001_11111111_11111111_11111111_11111011_01110111_01111100_11001100_11111111_11111111_11111111_11000010_01111101_01111100_11101100_11111111_11111111_11111111_10010100_01111110_01000111_11111100_11111111_11111111_11111111_00111100_01111101_10010100_11111111_11111111_11111111_11111101_01010101_01111101_10110111_11111111_11111111_11111111_11101101_01111100_01100000_11110101_11111111_11111111_11111111_11000110_01111100_10000010_11111111_11111111_01111011_10110100_11111111;
assign in[541] = 496'b01011100_11111111_11111111_11111111_11111111_01010000_01110011_11110010_11111111_11111111_11111111_11111111_01010000_01110111_11011011_11101101_10100011_01010100_11001011_01110111_01111100_01100100_01111100_01111100_01111100_00011011_01111101_01111101_01111110_01111101_01111101_01111101_01001100_01110001_11100100_11111001_11111001_00111010_01111100_01111100_01011010_11111111_11111111_11110001_01110001_01111001_01111100_10011111_11111111_11111111_11100010_00111111_01000000_01111100_11010100_11111111_11111111_11111111_11111111_11111111_11111111_11111111;
assign in[542] = 496'b11111111_11011010_10000011_00001001_11101111_11111111_11111111_00001110_01111000_00001101_01100010_11111111_11111111_11111110_01010110_10001011_11111111_11011111_11111111_11111111_11111011_01100111_00101010_10010000_01000110_11111111_11111111_11111111_10110100_01110100_01111110_01011101_11111111_11111111_11101010_11001101_00011001_01011110_11101000_11101000_00010010_01101110_01111110_10000011_11011001_11111111_01110001_01111110_01010111_10010000_11110100_11111111_11111111_10001001_11101110_11111110_11111111_11111111_11111111_11111111_11111111_11111111;
assign in[543] = 496'b11111111_11111111_11111111_10111000_10111101_01101011_00100010_00001110_01000001_01110100_01111010_00011110_01001000_01111101_01111110_01111101_01111101_01111101_11111111_11111111_10011001_01111101_01111100_01111100_01010011_11111111_11111111_01101101_01111110_01111101_01111101_01001101_11111111_11001101_01111100_01111101_01110101_00000100_11111011_11111111_00110101_01111101_01101110_11001101_11111111_11111111_11111111_01011000_01111100_10001110_11001000_11111111_11111111_11111111_01001001_01111100_01011110_01110101_10011011_01110010_01111101_01101011;
assign in[544] = 496'b11000000_01100101_01100101_01011101_11111111_11010110_01101110_10101011_11000110_10101000_11111111_11111111_00100000_00010110_11111111_11111111_11111111_11111111_11111111_01101010_11000011_11111111_11111111_11111111_11111111_11111111_01010001_10011001_11111111_11111111_11111111_11111111_11111111_10110011_01011110_00010011_00100110_10010110_11111111_11111111_11111111_10110101_01111011_10000100_10110110_11111111_11111111_11111111_00010110_00001101_11111111_11110101_11111111_11111111_11111111_10010011_01100111_00010111_01011110_11111100_10110111_10000001;
assign in[545] = 496'b11111111_10001000_01111100_01001000_11111111_11111111_11011001_00001100_01111100_01010111_11111111_11111111_11111111_11111010_01001101_01111101_00000110_11111111_11111111_11111111_10110110_01111101_01111100_11100000_11111111_11111111_11111111_10011110_01111110_01110001_11101100_11111111_11111111_11111111_00000001_01111101_00110011_11111111_11111111_11111111_11111111_00010001_01111101_10011111_11111111_11111111_11111111_11111111_00011001_01111110_10111010_11111111_11111111_11111111_11111111_01000011_01111101_11010101_11111111_01011011_01101010_11111111;
assign in[546] = 496'b11111111_11111111_11011000_01010111_01101011_11111111_11111111_11000010_01110110_01001100_11001110_11111111_11111111_10011100_01111001_00100111_11111111_11111111_11111111_10001011_01111000_00010100_11111101_11111111_11111111_11000100_01110110_00100110_11111010_11111111_11111111_11111111_01011011_01001011_11110000_11111111_11111111_11111111_11111111_01111101_00111001_10111110_11100010_11100010_11100010_11010111_00010001_01101001_01111101_01111101_01111101_01111101_01111101_11111111_11111111_11000101_10111100_10010111_10010000_11111111_11111111_11111111;
assign in[547] = 496'b10100111_11111111_11111111_11111011_11000011_01110011_01101000_11010110_00010000_01110001_01111101_11111111_01110100_01111101_01101000_01111101_00101101_10100110_11111111_00011011_01111101_01111101_01010111_11101101_11000000_11111111_00010101_01111101_01111101_01111101_01110000_01111010_11010000_01111100_01011100_11011101_11001011_10100010_10100110_10100010_01111101_10010101_11111111_11111111_11111111_11111111_10001000_01111101_10101111_11111111_11111111_11111111_11111111_10101100_01111101_01010010_00010100_01001100_10001011_01111101_01100010_00100010;
assign in[548] = 496'b11010000_01111111_00101111_11111111_11111111_11111111_00000000_01111111_10110000_11111111_11111111_11111111_11111111_01100000_01111111_11010000_11111111_11111111_11111111_11111111_01111111_01111111_00110000_01101111_00100000_11111111_10100000_01111111_01111111_01111111_01111111_01111111_11110000_01100000_01111111_00101111_10110000_01111111_01111111_11010000_01111111_01111111_00100000_01100000_01111111_00100000_11000000_01111111_01111111_01111111_01111111_00010000_11110000_11110000_01010000_01101111_00110000_11000000_11111111_11111111_11111111_11111111;
assign in[549] = 496'b11111111_11011110_01111101_11101010_11111111_11111111_11111111_10101110_01110001_11110001_11111111_11111111_11111111_11111111_00001000_00100011_11111111_11111111_11111111_11111111_11111101_01011111_10011100_11111111_11111111_11111111_11111111_11101011_01110101_10100110_11111111_11111111_11111111_11111111_11100101_01111101_10100110_11111111_11111111_11111111_11111111_10100101_01110111_11100100_11111111_11111111_11111111_11111111_10000100_01011100_11111111_11111111_11111111_11111111_11111111_10110011_01011100_11111111_11111111_11100010_10110000_11111111;
assign in[550] = 496'b00011111_01111101_10001000_11111111_11111111_11100010_01111000_01111101_11000001_11111111_11111111_11111111_11010010_01111100_01111101_11111111_11111111_11111111_11111011_01001001_01111100_01111101_01101010_01101010_01101010_11111001_01100011_01111011_01111000_01111001_01111011_01111101_10110101_01111100_00001101_11111111_11101011_01000000_01111010_00010111_01111100_11010000_11111111_10011100_01111100_00100000_01101011_01011101_11111101_11111111_01011000_01100101_11011011_01111100_10010110_11111111_11111111_10000100_11000101_11111111_11111111_11111111;
assign in[551] = 496'b11111111_10000010_01011001_11110101_11111111_11111111_10111101_01110010_11011000_11111111_11111111_11111111_11100011_01101000_10110011_11111111_11111111_11111111_11110001_01010100_10000101_11111111_11111111_11111111_11111111_00000111_00110101_11111111_11111111_11111111_11111111_11111111_01010100_11001001_11111111_11111111_11111111_11111111_11111111_00101001_00110010_11010101_11111111_11111111_11111111_11111111_11111100_10000111_01001100_01011110_00110001_00000101_00000101_11111111_11111111_11111111_11101111_11011101_10110110_11111111_11111111_11111111;
assign in[552] = 496'b10000010_10000010_10000010_10000010_10000010_01000101_01111101_01111101_01111101_01111101_01111101_10101100_01111101_01111101_00101001_11010110_10011110_10000001_00101000_01111101_01111101_11010110_11111111_11111111_11111111_01111101_01111101_00110111_11111111_11111111_11111111_11111111_01101111_01111101_00101001_11111111_11111111_11111111_11111111_00101001_01111101_01101111_11111111_11111111_11111111_11111111_10000010_01111101_01111101_10000010_11110010_11010111_11111111_11010110_01111101_01111101_01111101_01100001_01111101_01111101_01111101_01100001;
assign in[553] = 496'b00110101_11111111_11111111_11111111_11111111_11000100_01111101_11101101_11111111_11111111_11111111_11111111_11011100_01111101_10100011_11000101_10101110_11110000_11111111_11011100_01111101_01111010_01000111_01100110_01000011_11111111_11011100_01111110_10100100_11111111_00010001_01011010_11111111_10101101_01111101_11011001_11111111_00010101_00110101_11111111_10000011_00111001_11111110_11100001_01110101_11000011_11111111_00110010_00010100_11101100_00111100_00101010_11111100_11111111_11001101_01110101_01110101_01101011_11010011_10111000_10011110_11101101;
assign in[554] = 496'b11011010_01001001_11111111_11111111_11111111_11111111_10100010_00101011_11111111_11111111_11111111_11111111_11111111_00010101_10001011_11111111_11111111_11111111_11111111_11111111_01010100_10101010_11110111_11010010_11111011_11111111_11111111_01110101_11010111_00101000_01111110_01010100_11111111_11111111_01101101_00110111_00001110_00001010_01010110_11111111_11111111_01110101_01101000_11011101_00111011_10100101_11111111_11111111_01000100_01111001_01110111_10001111_11111110_11111111_11111111_11111111_10011100_11010001_11111111_11111111_11111111_11111111;
assign in[555] = 496'b11100010_10100111_01001011_01101010_01111101_01000111_01111101_01111101_01111101_01101001_00011000_01101010_00011110_01111101_01111101_00100000_11111101_11111111_11111111_11010011_01111101_01011110_11111101_11111111_11111111_11111001_01010001_01111011_11100101_11111111_11111111_11111111_11101011_01111101_00100100_11111111_11111111_11111111_11111111_11101011_01111101_10110001_11111111_11111111_11011001_11111011_11101011_01111101_00101111_11001000_10101110_01110000_01101001_11111110_10011010_01111101_01111101_01111101_01111101_10111001_10000001_10000001;
assign in[556] = 496'b11001110_01001100_01111101_01111100_01111100_11001000_01011010_01111100_00001010_11101100_10010101_11110001_01100110_01111011_10000110_11111111_11111111_11111111_10101101_01111100_00011111_11111111_11111111_11111111_11111111_10011111_01111101_00110000_10000010_00110001_00110101_11000101_11110011_01010110_01111100_01111100_01111101_01111100_00011001_11111111_00011000_01111100_00111101_00011001_00011001_10110101_11111111_01101000_01111100_00101001_10011000_10111100_10011000_11111111_00101110_01111000_01111100_01111101_01111011_11101100_10001110_10010001;
assign in[557] = 496'b10010110_01111101_11001111_11111111_11111111_11111111_01001010_01101011_11110011_11111111_11111111_11111111_11010110_01111000_00010101_11111111_11111111_11101010_11111111_10000101_01111101_10111111_11111111_11111111_01000010_11111111_01010000_01011101_11111110_11111111_11010101_01111011_11101010_01111010_00110010_11111111_11111111_00001100_01111101_00001111_01111101_01111101_00001100_11101100_01010000_01011111_00110111_00111011_00110101_01111101_01111100_01110111_10101001_11110011_11111110_11111101_10101000_10000001_11010011_11111111_11111111_11111111;
assign in[558] = 496'b11111111_11010001_00110000_01010000_11000000_11111111_11111111_01010000_01111111_01111111_01111111_11111111_11111111_10100000_01111111_10110000_01000000_01111111_11111111_11111111_00110000_01111111_01010000_01111111_00010000_11111111_11110000_01111111_01111111_01111111_10100000_11111111_11111111_00010000_01111111_01010000_11010000_11111111_11111111_01000000_01101111_01111111_00000000_11111111_11111111_11111111_11000000_11000000_01111111_00101111_11111111_11111111_11111111_11111111_11111111_01010000_01111111_11110000_11111111_10010001_01111111_11100000;
assign in[559] = 496'b10001000_11000100_11111001_11111111_11111111_00011011_01010000_01110101_01100101_10100101_11111111_10110011_11111111_11111111_11101011_10001110_01101111_10011011_00001000_11111111_11111111_11111111_11111111_10010101_01111000_01110011_10110011_11111111_11111111_11111111_11111110_01001000_10110101_01011100_00001001_11111111_11111111_11110000_01000010_11111111_11011000_01000100_01101111_01010110_01110100_01111110_11111111_11111111_11111110_11010110_10110000_00110100_01101000_11111111_11111111_11111111_11111111_10110101_01111000_11101011_10001000_01101100;
assign in[560] = 496'b11111001_10011010_10000001_00000000_11100101_10100010_01011011_01111011_01110110_01110111_01111110_00101110_01111001_10001000_11011110_11111111_11110111_10110000_01111110_00010110_11111111_11111111_11111111_11111111_11111111_00111001_01001100_11101110_11111111_11111111_11111111_11111111_10111010_01101100_01110011_00010001_11010111_11011110_11110101_11111111_11010110_00010100_01111001_01111110_01111110_10101111_11111111_11111111_11111111_00101100_01111000_10001100_11111001_11111111_11111111_11101001_01111100_00000100_11111111_11111111_00111101_01111001;
assign in[561] = 496'b01111011_01111100_01010100_10011101_00100001_01111100_01110100_10000110_11101100_11111111_11110100_01001110_01100110_10111010_11111111_11111111_11111111_11001100_01111011_00001110_11111111_11111111_11111111_11111111_00010001_01111100_10110111_11111111_11111111_11111111_11101101_01101011_01111011_01011111_11100111_11110001_11110110_00001111_01101011_01100000_01111100_01111011_01111100_01010000_01111011_00100001_10110000_01110101_01111100_01111101_01111100_00010100_11110111_11111111_11100110_00110100_01111100_01011011_11111000_10001011_01100100_10101100;
assign in[562] = 496'b11111110_01011110_10100000_11111111_11111111_11111111_11111001_01111110_10011101_11111111_11111111_11111111_11111111_11111001_01111110_11000010_11111101_11011001_11111111_11111111_11100011_01111110_10010000_01011000_01111111_11111111_11111111_11000100_01111110_01111110_01000101_10010110_11111111_11111111_10110001_01111110_00100110_11111111_11111111_11111111_11111111_00011111_01110110_11011110_11111111_11111111_11111111_11110111_01110100_01001000_11111111_11111111_11111111_11111111_11110011_01111110_10001000_11111111_11111111_10100111_11101000_11111111;
assign in[563] = 496'b11111000_01010110_01111000_10111100_11111111_11111111_00010001_01111101_00110111_11111111_11111111_11111111_11100100_01011100_01101000_11101011_11111111_11111111_11111111_10001010_01111101_10001111_11111111_11111111_11111111_11111111_01000111_01101001_11101111_11111111_11111111_10001110_11010100_01111011_10010001_11111111_11111001_00000110_01110101_10111000_01111011_11010001_11010100_01011000_01111001_10010000_10001011_01110100_01001001_01111000_01011100_11000010_11111111_10111101_01101101_01110100_00001011_11101010_11111111_11111111_11111111_11111111;
assign in[564] = 496'b11111111_11111111_11111111_11111010_10100011_11100101_11111111_11111111_11110110_01000000_01111110_00111001_01101011_01011010_00000000_01001011_01111110_01111100_11111111_11111001_10000010_01111110_01111110_01110100_10011100_11111111_11111111_10010111_00100110_11000110_11110010_11111111_11111111_11110111_01100100_11100000_11111111_11111111_11111111_11111111_10001111_00100111_11111111_11111111_11111111_11010010_11111111_00001110_10001100_11111111_11111100_00101000_00110101_11111111_00001110_10010001_11101111_00110001_01001001_01011111_01001010_10011101;
assign in[565] = 496'b11111111_10011101_00100111_11111111_11111111_11111111_11111111_00101111_10101010_11111111_11111111_11111111_11111111_11111010_01011110_11111000_11111111_11111111_11111111_11111111_10110100_00100101_11111100_11111110_11111111_11111111_11111111_00110010_00001110_01010110_01000101_11111111_11111111_11011110_01111000_01011001_00010011_00100110_11111111_11111111_00010100_00110101_11010001_01001010_11011101_11111111_11111111_01100001_00010111_01001011_11011110_11111111_11111111_11111111_10100010_10011111_11110110_11111111_11111111_11111111_11111111_11111111;
assign in[566] = 496'b11111011_11111111_11111111_11111111_11111111_01011010_11111111_11111111_11111111_11111111_11111111_11010111_01100010_11111101_11111111_11111111_11111111_11111111_11110000_01111000_11011100_10111001_00010100_00011001_10100010_11111111_01110100_01001000_01111110_01110010_01111001_01111111_11111111_01110100_01011100_10010001_11110101_11110111_01001100_11111111_00110101_00101101_11000101_11011111_10000111_01110100_11111111_11011001_01011111_01111100_01111110_01111101_10010100_11111111_11111111_11111111_11010000_10100110_11001000_11111111_11111111_11111111;
assign in[567] = 496'b00101010_01110110_00111000_01101110_00001011_10000011_01101001_11100011_11111111_11111010_01110010_11111100_01100100_10110100_11111111_11111111_11111111_10110000_11000100_01111000_11101001_11111111_11111111_11111111_11111111_11000101_01110011_11111001_11111111_11111111_11111111_11111111_11111100_01011010_00000000_11111111_11111111_11111111_11111111_11111111_11001001_01101000_00110101_00001110_11100100_11001110_11111111_11111111_10000001_01110110_00010100_11101001_10100101_11111111_11111000_01101110_01100100_01000010_01101111_10111111_10000001_10001011;
assign in[568] = 496'b11111111_11111011_00011101_01111000_01111110_11111111_11111111_00001001_01111000_00001001_11011100_11111111_11111111_11110001_01111000_10100000_11111111_11111111_11111111_11111111_10101010_01111101_10110100_11111111_11111111_11111111_11111111_11100111_01111101_01110011_11111111_11111111_11111111_11100111_01000001_01101001_10111001_11111111_11111111_11011000_01011111_00110010_11100111_11111011_11111111_11111111_01010000_00001001_11001001_10000010_01011111_11001101_11111111_01111110_01101110_01110011_00011110_10110100_11111111_11110001_11111111_11111111;
assign in[569] = 496'b10000100_01101100_01111101_00111011_11101101_01001010_01101001_00000101_10010100_01101000_00011111_01000110_00111110_11100101_11111111_11111111_00000111_01110001_01010010_11111010_11111111_11111111_11111111_10100011_01111000_10100110_11111111_11111111_11111111_11111111_10100011_01110111_11100101_11111111_11111111_11111111_11111111_00001110_01110001_00101000_11100101_11101011_11011000_10111100_01011001_01000011_01100110_01110101_01110001_01111000_01111100_01111101_10100110_11110001_11011000_11011000_11100000_01011011_01011001_11111111_11111111_00100011;
assign in[570] = 496'b11111111_11111010_10110000_00001011_10001000_11111111_11101001_01010100_01111110_01110110_01011100_11111111_11111111_00100010_01111101_10000011_11110101_11111111_11111111_11111111_00110110_01001010_11111100_11111111_11111111_11111111_11111111_11011101_01010101_00010111_11110001_11111111_11111111_11111111_11111111_11100000_01100011_10011000_11111111_00001101_01000011_01100011_01110110_01100101_11000011_11111111_01110011_01110110_01100011_10001000_10011011_11011010_11111111_11101010_11110111_11111001_11111111_11111111_11111111_11111111_11111111_11111111;
assign in[571] = 496'b10011110_01111110_01110011_11101010_11111111_11100110_01011100_01111110_00001010_11111111_11111111_11111111_10001100_01111110_01101010_11110001_11111111_11111111_11111011_01110110_01111110_10100100_11111111_11111111_11101010_10101100_01111110_00101111_11111011_11111111_11010001_01110000_00000010_01111111_10010000_11111111_11111011_00111010_01111110_11100011_01110100_00111110_00101001_01101110_01111110_01101100_11111111_11000000_01011001_01111110_01011101_01001111_10101010_11111111_11111111_11111010_10100000_00001000_10010010_11111111_11111111_11111111;
assign in[572] = 496'b11010110_00111001_01111101_01111101_01111101_11000110_01101000_01111101_01110111_00110110_01111001_11011011_01110101_01111101_01110010_11000111_11111111_00111011_01000101_01111101_01110100_10110101_11111111_11111111_01010101_01111101_01110010_10101110_11111111_11111111_11000100_01111000_01111101_00101011_11111111_11111111_11100110_01001011_01111101_01111101_00001100_10000001_01101000_01010010_01111101_01110100_01111101_01100100_01011011_01111101_01111101_01110100_11011001_00011101_01111101_01111101_01111101_01111101_10100111_10100110_10001001_11000010;
assign in[573] = 496'b11111111_00010011_01111101_01100000_00000110_11111111_10101101_01111101_00101011_11110010_11111101_11111111_11111111_01001001_01010101_11110101_11111111_11111111_11111111_11111111_00111011_10001010_11111111_11111111_11111111_11111111_11001010_01010110_01110000_11101000_11111111_11001000_10000001_01111110_01100111_00010101_11101110_00011010_01111110_01111011_00001001_11100110_11100011_00110011_01111110_01000001_01111010_00000011_00011000_01101100_01111110_00111010_11011110_00001001_01110001_01101010_01000101_10100000_11111011_11111111_11111111_11111111;
assign in[574] = 496'b10011101_00110101_01001111_01101101_00001001_01010001_01110000_00110100_00011010_10000100_00111100_00011011_00111111_11011010_11111111_11111111_11111111_11111111_01011010_11000110_11111111_11111111_11111111_11111111_11110101_10001010_00110111_10011010_11001000_11001100_11110000_11111111_11110011_10110101_00111010_01111001_01111101_10000100_11111111_11111111_11111111_11110011_01010010_01101010_10110101_11111111_11111111_11111111_00101001_01101111_10011001_01000100_11011110_11111111_11100010_01110111_01111010_01111001_00100011_01101101_00011000_11010010;
assign in[575] = 496'b11111111_11111111_11111111_11111111_11111111_00011111_01110000_01110001_01110010_00111101_11000110_10110011_11000011_10010101_00111011_10001011_00101011_01001101_11111111_11111111_11111111_11110101_00011100_10101101_01110001_11111111_11111111_11111111_11111111_00011100_10110001_00110100_11111111_11111111_11111111_10011001_01001001_11111000_00010010_10100011_10101100_00110001_01011010_11001111_11111111_00101110_00001001_10010100_10110010_11111111_11111111_11111111_01011111_11111111_11111111_11111111_11111111_11111111_11110000_11111111_11111111_11111111;
assign in[576] = 496'b11111111_11111111_11111111_11111101_11100010_11111111_11111111_11111111_11110111_00101111_01111110_10101010_10101000_10000010_00001010_01011011_01111110_01111110_01000101_01010100_01111100_01111110_01110010_01000100_10100011_11111111_11000100_01101100_01100001_11010011_11111111_11111111_11111111_01011101_01100010_11010011_11111111_10100011_10011110_10111011_01110000_11000000_11111111_10100000_01111100_00111010_10000100_00001110_11111111_10111101_01110001_00110111_11101000_10001010_00110001_00010101_01011111_00000011_11111000_00101111_11011100_11111111;
assign in[577] = 496'b11111111_11111111_10100101_01111110_10101100_11111111_11111111_11010111_01110011_00001001_11111111_11111111_11111111_11111011_01000001_01000101_11111011_11111111_11111111_11111111_00000101_01100001_11110100_11111111_11111111_11111111_11101100_01110000_10011101_11111111_10100101_11001011_11111111_10011010_00111010_11111111_10110011_01111110_10111000_11111111_00100110_10100011_11101001_01101100_10000111_11111111_11111111_00011011_00100001_01001000_01000000_11111111_11111111_11111111_11010011_01101001_01000000_11010111_11111111_11111111_11111111_11111111;
assign in[578] = 496'b11111011_10110101_10100000_11110101_11111111_11000101_01001010_01111110_01111110_01011100_11100101_11101011_01100010_01010101_01111110_00000011_01101110_00100010_10001011_01100001_11110111_01111110_11001001_00010111_00101001_00001010_00101110_11010010_01100000_11110110_00001111_00101001_10001011_01011001_00111011_10000110_11101111_01110000_10101010_11010111_01011110_01001100_11111111_00101111_01010101_11111011_11111111_11111101_11111101_10101001_01111000_10111111_11111111_11111111_11111111_11111110_01110111_10000010_11111111_10011000_00111010_11111100;
assign in[579] = 496'b01001001_00000101_01101100_10010111_11111111_01110000_11011110_11111111_11100010_11101101_11111111_10110111_00110010_11111111_11111111_11111111_11111111_11111111_11110011_01100100_11100110_11111111_11111111_11111111_11111111_11111111_10010101_01010000_11011110_11111111_11111111_11111111_11111111_11111111_10100110_01011101_01000100_11101100_11111111_11111111_11111111_11110110_00110110_00100010_11111000_11111111_11111111_11111111_10011000_01001011_11111111_11111111_11111111_11111111_11111111_11100010_01011100_00101011_10000111_11111111_11101100_10010101;
assign in[580] = 496'b00111000_11111111_11111111_11111111_11111111_01011101_01000010_11111111_11010110_11110100_11111111_11111111_00000010_01111110_11010011_00110100_10000001_11111111_11111111_10010000_01111110_00100001_01110001_00000010_11111111_11111111_10010000_01111110_00110110_01111010_00000010_11111111_11111111_11011110_01111100_10110101_00101011_00101010_11111111_11111111_11111111_01111001_10010101_11010011_01111101_11011000_11111111_11111111_01100011_10110001_11111111_01001000_10101000_11111111_11111111_11000000_11011100_11111111_10001111_11111111_11111111_11111111;
assign in[581] = 496'b11111111_11111111_11111111_10110001_01110010_11111111_11111111_11111111_11111101_00110010_01110000_11111111_11111111_11111111_11111111_00001011_01111100_00010101_11111111_11111111_11111111_10111101_01111010_00111101_11111001_11111111_11111111_11010111_01110011_00111101_11110000_11111111_11111111_11101000_01001000_01100101_11001010_11111111_11111111_11111110_00010111_01111011_10101000_11111111_11111111_11111111_10101010_01111101_10001101_11111111_11111111_11111111_11111111_01000000_01001101_11111011_11111111_11111111_11111111_11111111_11111111_11111111;
assign in[582] = 496'b11111111_11111111_11111111_11111111_11110000_11111111_11111111_11111111_11111111_11110000_01010000_11111111_11111111_11111111_11111111_11000000_01100000_01111111_11111111_11111111_11111111_10110000_01111111_01111111_00000000_11111111_11111111_10100000_01111111_01111111_11100000_11111111_11111111_11000000_01101111_01111111_10110000_11111111_11111111_11000000_01101111_01101111_11010000_11111111_11111111_11111111_01100000_01111111_10110000_11111111_11111111_11111111_11111111_01111111_00000000_11111111_11111111_11111111_11111111_11111111_11111111_11111111;
assign in[583] = 496'b11111111_10110101_01001001_00011011_01000110_11111111_11010000_01110011_11100001_11111111_11111111_11111111_11111111_00000011_00100011_11111111_11111111_11111111_11111111_11111111_10000110_01010010_10100001_10111010_11001111_11111111_11111111_11111100_10001011_00011011_00111101_01100001_11111111_11111111_11111111_11111111_11111111_10001100_00011101_11111111_11100001_11101110_11011011_10101011_01010110_11010100_10101000_01011101_01110101_01100111_01100011_00001001_11111111_01111100_00110010_10000101_11101100_11111111_11111111_11111111_11111111_11111111;
assign in[584] = 496'b11001010_00101011_01111001_01111101_01010011_00110010_01111101_01111101_01011101_01101101_01111101_01010011_01111100_10000101_11011111_11111110_11110100_01010101_01111101_10001011_11111111_11111111_11111111_11111111_01010001_01011010_11111101_11111111_11111111_11111111_11111111_01010110_00101011_11111111_11111111_11111111_11111111_11000001_01111101_00010111_11111111_11111111_11111111_10010000_01101001_01111101_01010100_11110110_10111111_01001000_01111001_01111101_01010011_01111101_01010111_01111101_01111101_01111101_00101111_01111110_01001100_10011011;
assign in[585] = 496'b01111100_11010110_11111111_11111111_11111111_10111111_01110111_11110000_11111111_11111111_11111111_11111111_00010010_01001001_11111111_11111111_11111111_11111111_11111111_00110011_00101100_11111111_11101110_10111001_11010100_11111111_00111111_01000101_01001010_01110100_01111101_01110011_11111111_01010110_00111001_10101011_10111111_10110101_01111101_11101101_01110110_11000010_11111111_11111111_00011111_01010110_11100001_01111101_11100000_11111111_11111111_00111101_10010101_11111111_10001001_11110010_11111111_11111111_01011111_11111111_11111111_11100100;
assign in[586] = 496'b11111111_11111111_10111011_10101001_11111111_11110111_10010100_00111011_01111000_01111100_11110100_11110110_01010000_01011000_00001011_01111000_01001001_11111111_11110100_01100000_01111101_01100100_01110001_00001111_11111111_11111111_11111100_11011000_11011110_00001110_10000111_11111111_11111111_11111111_11111111_11111111_00111110_10110000_11111111_11111111_11111111_11111111_11101000_01101110_11011010_11111111_11111111_11111111_11111111_10001000_00101001_11111111_11111111_11111111_11111111_11001010_01100001_11000111_11111111_01101010_10100101_11111111;
assign in[587] = 496'b11111111_00000010_01111110_01001101_11101100_11111111_11111111_00010101_00111100_00011011_00010000_11111111_11111111_11111111_10100100_01000001_11000111_01000111_11111111_11111111_11111111_11010101_01111011_01110000_00100100_11111111_11111111_11000000_01000100_01111110_00011001_11110011_11100000_00110101_01111000_00101000_01100010_10100011_11111111_01011000_00111110_11011000_11111111_01000100_10100000_11111111_00111001_11111011_10101111_11111111_01000100_10100110_11111111_11011000_11111111_00001101_01000100_01100100_11011011_11101011_10001111_11011110;
assign in[588] = 496'b11111111_11111111_11111111_11111111_11111111_01010101_01111111_01111111_01011100_00010101_11101011_01011100_10100100_00001110_01101010_10011101_01010101_01000000_11001000_11101011_01000111_01000000_11111111_10110010_01111111_00111000_01110001_01010101_11011101_11111111_10101011_01111111_10001111_10111001_11111111_11111111_11111111_10001111_01110001_11111111_11111111_11111111_11111111_11111001_01100011_10001000_11111111_11111111_11111111_11111111_10010110_01101010_11110010_11111111_11111111_11111111_11110010_01101010_00000111_11111111_00010101_01001110;
assign in[589] = 496'b11111111_11110100_01101110_10100101_11111111_11111111_11111111_10111010_01111011_11011001_11111111_11111111_11111111_11111111_00100001_00111101_11111111_11111111_11101101_10011000_00000011_01111101_00010111_11101001_11111111_10011000_00010011_01111010_01010110_01001000_01110101_10101110_11111111_11010010_01101101_11101000_11111111_00111100_10001000_11111111_00010010_00001010_11111111_11111011_01100110_11001011_11111111_01100000_11001110_11111111_10110110_01001010_11111101_11011100_01010010_11111100_11111111_11010111_11100101_11111111_11111111_11111111;
assign in[590] = 496'b00100011_11111111_11111111_11111111_11111111_11111111_01010000_11111111_11111111_11111111_11111111_11111111_11111111_01000010_11111111_11111111_11111111_11111111_11110111_10001011_01100110_00111001_00100101_10011001_11101101_11011011_10011001_00001011_11111111_11100001_00001100_01011000_11111111_10101101_10001111_11111111_11111111_11111111_11000100_11111111_10011110_10101001_11111111_11111111_11111111_11111111_11111111_10001000_11000000_11111111_11111111_11111111_11111111_11111111_00010000_11011101_11111111_11111111_11111111_11110110_11111111_11111111;
assign in[591] = 496'b11111111_11111111_11111111_11111111_11111111_01101111_11111000_11111111_11111111_11111111_11111111_11001111_01111011_11001011_11111111_11111111_11111111_11111111_11111111_00100101_10001010_11100100_10101100_10011011_10110101_11111111_10000111_01011011_01100010_00100111_00011000_00110010_11111111_10111010_01100100_11101101_11111111_11111111_11001100_11111111_11000011_01010100_11111111_11111111_11111111_10100000_11111111_11000101_01110101_11111101_11111111_11111111_11111110_11111111_11101001_01101111_11111101_11111111_11111111_01011000_11111100_11111111;
assign in[592] = 496'b10100000_10100000_00011000_11111101_11111111_10100010_11111111_11111111_11111111_11111111_11111111_01111101_00000111_11111111_11111111_11111111_11111111_11111111_01010110_01101110_10001001_11010101_11010101_11010101_11101111_11100001_00101100_01111101_01111101_01111101_01111101_00101101_11111111_11111100_00000100_01111101_01111101_01101101_10010011_11111111_11111111_10100010_01111101_01111101_10011001_11111010_11111111_11111111_11111101_10011001_01111000_01111101_00111100_11111111_11111111_11111111_11111111_11100110_00100000_11111111_11111111_11111111;
assign in[593] = 496'b11101010_10001010_10001010_11111001_11111111_11111011_01000011_01100100_01101110_10010000_11111111_11111111_10110100_01111000_11011110_10001101_00101010_11111111_11111111_10001010_01110011_11111111_00111101_00000000_11111111_11111111_11001011_01110111_00111110_01111011_01001011_10111011_11111111_11111111_10111101_00101110_01001011_11110110_11111111_11111111_11111111_11101110_01001101_11001101_11111111_11111111_11111111_11111111_00101001_00101000_11111111_11111111_11111111_11111111_11001101_01111010_11000111_11111111_11111111_01111010_10110111_11111111;
assign in[594] = 496'b00010001_01101001_01111110_01111110_01111110_01010100_01111101_00110000_00001101_10100011_01011111_00110011_01110010_10101000_11111111_11111111_11111111_00001110_01100010_00010010_11111111_11111111_11111000_11101110_01011001_01111110_11000100_11111111_11111111_00000110_01110110_01111110_01100111_11110100_11111111_11111111_10111100_01111100_01101100_00101111_11111111_11111111_11101110_01001101_01111110_10000100_01010000_10100101_10000010_01110100_01111110_01001000_11110111_01101011_01111110_01111110_01111001_00011011_11110110_11001100_11111000_11111111;
assign in[595] = 496'b11111111_11111111_11111111_11111111_11111111_11000110_00110101_01111110_01111110_01100100_10111000_10101011_01101110_00010111_01010101_01011011_01000000_01110010_01001010_10110111_11101111_01011000_00101101_10101110_01111110_01110110_10010100_01010101_01101111_11010111_00010101_01111110_01110111_01110111_10000111_11100100_11111111_00111110_00101100_11111111_11111111_11111111_11111111_10101011_01111110_10110100_11111111_11111111_11111111_11111111_01000011_01000010_11111110_11111111_11111111_11111111_11010100_01111011_10100111_11111111_10010001_01011011;
assign in[596] = 496'b11111111_11111001_01101010_11000000_11111111_11111111_11111111_11010101_01111111_11100100_11111111_11111111_11111111_11111111_00000111_01010101_11111111_11111111_11111111_11111111_11111111_01000000_00010101_11111111_11111111_11111111_11111111_11101011_01111111_10101011_11111111_11111111_11111111_11111111_11010101_01111111_11110010_11111111_11111111_11111111_11111111_11010101_01111111_11101011_11111111_11111111_11111111_11111111_11010101_01111111_11101011_11111111_11111111_11111111_11111111_11001110_01111111_11111111_11111111_11011101_01110001_11110010;
assign in[597] = 496'b01011101_11100001_11111111_11111111_11111111_11111011_01011001_11111111_11111111_11111111_11111111_11111111_10110110_00110001_11111111_11111111_11111111_11111111_11111111_10011010_00001111_11111111_11111111_11111111_11111111_11111111_00011000_10011100_11111111_11111111_11111111_11111111_11111111_01010001_11100001_11111111_11111111_11111111_11111111_11101100_01011001_11110011_11001111_10101100_10010010_00001100_11010011_00100110_00100110_00010001_10011010_10110100_11011011_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111;
assign in[598] = 496'b11111111_10010110_01000001_11111111_11111111_11111111_11110000_01100011_10001111_11111111_11111111_11111111_11111110_00011111_01100101_11100111_11111111_11111111_11111111_10100100_01111100_10011010_11111111_11111111_11111111_11111111_01000011_00110111_11111111_11111111_11111111_11111111_10110001_01110111_11011000_11111111_11111111_11111111_11111111_01001110_01100000_00000110_00000110_00000110_00000110_00101100_00111110_00100011_00011111_00101001_00101001_00100110_10000011_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111;
assign in[599] = 496'b10000010_10000010_10000010_10111100_11111111_10001011_11000101_11001111_10100111_01001111_10001110_01000000_11111111_11111111_11111111_11111111_11101010_01110010_01000100_00010011_11010000_11111100_11110001_00110001_01000101_11101100_10011100_00010100_00101100_00010101_10101101_01001000_11111111_11111111_11111111_11111111_11111111_11100111_01011000_11111111_11111111_11111111_11111111_11111111_00101010_10010010_11111111_11111111_11111111_11111111_10011110_01000110_11111101_11111111_11111111_11111111_10100001_01000000_11100010_00011010_01001110_11100010;
assign in[600] = 496'b11111111_11111111_00010000_10001110_11111111_11111111_11111111_11100101_01100001_11101111_11111111_11111111_11111111_11111111_00010111_00000110_11111111_11111111_10101010_00110110_01010100_01111100_10001100_11111011_11111111_11001011_11010010_01110110_01001100_01011111_01100110_11011010_11111111_10011100_01001100_11111101_11111111_00101101_10010100_11111111_01010001_10011101_11111111_11111111_00100011_10000010_11001011_01011001_11111011_11111111_11011101_01101110_11101010_00011111_10100010_11111111_11111111_10011100_10011110_11111111_11111111_11111011;
assign in[601] = 496'b11001111_10101110_10001000_10001000_10111010_10001111_01111000_01010011_01010011_01010011_01111000_11010111_01111010_10100101_11111111_11111111_11111111_11100111_11001000_01111100_11100100_11111111_11111111_11111111_11111111_11110001_01101010_00100110_11101010_11111111_11111111_11111111_11111111_11010110_00101110_01010011_00001000_10101011_11010110_11111111_11111111_11111111_11011011_01011000_01100110_00011110_11111111_11111111_11101010_01011101_10001100_11110111_11111111_11111111_11111111_00010110_00010010_11111111_11111001_10100101_01011111_00001110;
assign in[602] = 496'b11011010_10000100_00100011_00101101_10100111_00011101_01101101_01001000_00110011_01100100_01111101_01110111_01000001_11000100_11111111_11111111_11011100_01111100_00101011_11111110_11111111_11111111_11111111_11111111_10101101_11010010_11111111_11111111_11111111_11111111_11111111_10011111_11111111_11111111_11111111_11111111_11111111_11111000_01010111_11111111_11111111_11111111_11111111_11111011_01000011_01111101_11101111_11111111_11100010_10101010_01000110_01111100_10000111_00001011_01010111_01111011_01111101_01111000_10010001_10010100_10111001_11100101;
assign in[603] = 496'b11000001_01011100_01011111_00001111_00000100_10111111_01101101_10001010_11111001_11111111_11111111_11111111_01000010_10100000_11111111_11111111_11111111_11111111_11111000_01111000_11001011_11111111_11111111_11111111_11111111_11111111_10110000_01011001_01011011_01000100_11000111_11111111_11111111_11111010_01011110_00100010_00100000_00110100_11111111_11111111_10111001_01101000_11111111_11111111_11111111_11111111_11111111_10100100_01101101_11111000_11111111_11111111_11101010_11111111_11111010_01001110_01100000_01101100_01100101_11111001_10101001_10000001;
assign in[604] = 496'b01101000_01110010_01110011_01010011_11011010_00100000_11011010_11111111_11111101_10100101_01101011_01011011_11101101_11111111_11111111_11111111_11111111_10010001_10010011_11111111_11111111_11111111_11111111_11111111_11110010_11010011_11111111_11111111_11111111_11111111_11111111_11111111_10110110_11111111_11111111_11111111_11111111_11111111_11010100_10000101_11111111_11111111_11111111_11111111_11111111_00101011_01101001_11011100_11111111_11111100_10011110_11001110_01100010_00000100_01100100_10001010_11101100_00010010_01010001_11010110_11111100_01011110;
assign in[605] = 496'b11010101_10001000_11001110_11011010_11111111_10010111_01111011_01111110_01111110_01111000_10010100_11011100_01010111_10101101_11111100_11111100_11101011_11001001_10100000_00100110_11111111_11111111_11111111_11111111_11111111_11001011_01111001_10111010_11111111_11111111_11111111_11111111_11111111_10010100_01101100_01110000_00100110_10000100_11000100_11111111_11111111_11011011_00001100_00011001_01111001_00101110_11111111_11111111_11111111_11111111_11010010_01110111_10001100_11111111_11111111_11111111_11110111_01100000_01000010_11111111_01011100_01010110;
assign in[606] = 496'b11110111_10100101_11111111_11111111_11111111_11111111_10101111_01111100_10001110_11101100_11101100_11111111_11111111_11111001_00101011_01111110_01110001_01110010_11111111_11111111_11111111_11001000_01111101_01111100_01100110_11111111_11111111_10100001_01101001_01111010_00111000_11101000_11111111_10000011_01111101_01100111_10110001_11111111_11111111_11111101_01010111_01100001_11011011_11111111_11111111_11111111_11100101_01111110_00011001_11111111_11111111_11111111_11111111_11111111_01000111_01000110_11111100_11111111_11111111_01111001_00011001_11111111;
assign in[607] = 496'b11111111_11111111_11111111_11111111_11111111_01110001_11100010_11111111_11111111_11111111_11111111_00010010_01111100_10010001_11000011_10111100_11011011_11111001_01111011_01111101_01111101_01111110_01111101_01101111_01011010_11101000_01111001_01010110_11111111_11110110_11011011_01101101_11111111_01000111_01010110_11111111_11111111_11100101_01101110_11111111_00101010_01010110_11111111_11111111_00001001_01111100_11111111_00101010_01100010_11111011_10110110_01111001_00111010_11111111_11010001_00000100_11110111_00110010_01011111_11111111_11111111_11111111;
assign in[608] = 496'b11111111_11111111_11101101_01010100_10000001_11111111_11111111_11101100_01001110_00011110_11111111_11111111_11111111_11110001_01000001_00100100_11110111_11111111_00100011_01011110_01110111_01001100_11111010_11111111_11111111_10111100_10010010_01101111_11101001_11111111_11111111_11111111_11111111_00111010_00010011_11111111_11111111_11111111_11111111_11110101_01110011_11101101_11111111_11111111_11111111_11111111_11101110_01101101_10001001_10100100_10100100_10001010_10011011_11111111_10110010_00010000_00001100_00001001_10011100_11111111_11111111_11111111;
assign in[609] = 496'b11111111_11111111_11111111_11111111_11111111_10001100_10000001_10100001_11001110_11111111_11111111_01111101_01111101_01111110_01111101_01111100_00110100_11100010_10010010_11001011_11001011_11001011_01100001_01111101_01011010_01111011_01111101_01111110_01111101_01111101_01110011_01111101_11010110_11010001_11010001_11010001_11010001_11101010_01011101_11111111_11111111_11111111_11111111_11111111_11101100_01110100_11111111_11111111_11111111_11111111_11111111_10111100_01111101_11111111_11111111_11111111_11111111_11111111_01001100_11111111_11111111_10011111;
assign in[610] = 496'b10111011_00101001_01111000_01111110_01110011_00110110_01110100_00010111_10101110_10111111_10100000_10010101_01101000_11100010_11111111_11111111_11111111_11111111_00001110_00010001_11111111_11111111_11111111_11111111_11111111_10011010_01100000_11000111_11111111_11111111_11101001_11111111_11111111_00000100_01110101_01100111_01111000_01010001_11111111_11111111_11111111_00111001_01101100_10011111_11011001_11111111_11111111_10111001_01111101_10101011_11111111_11111111_11111111_11111111_10010011_01101000_10101101_11001100_11001100_00111100_01001010_01100010;
assign in[611] = 496'b11111111_11111100_11011011_10110110_11110011_11110101_10000100_01011111_01110111_01111001_01110100_11101011_01010110_01100001_01011110_10101011_10111101_01111001_01000111_01011011_11100111_11111111_11111111_11111111_01101111_01111110_10010100_11111111_11111111_11111111_11011000_01111101_01111111_11000111_11111111_11111111_11100101_00110010_01111110_01110100_00110010_11111111_11101000_11011011_01110100_00100111_10010000_01110011_01010100_01111000_01110111_00111111_11110101_11111111_11110110_10011111_01011000_01010111_11011111_11111111_11111111_11111111;
assign in[612] = 496'b10010101_00110110_01100101_01111101_11010110_00111101_01111000_00111000_00101001_01101111_01001011_10111010_01111101_11000101_11111111_11100011_01101000_00100001_10111110_01111100_00000011_11100101_00101101_01110101_11101001_11111111_00010000_01001110_01111110_01111101_10010111_11111111_11111111_11100010_01100001_01110100_01101110_01101001_11110101_11111111_00101010_01000010_11011010_10101010_01111101_10111110_10010111_01011101_11111010_11110100_00101011_01101110_11111111_01010010_01010011_01101110_01110010_01100010_11001011_00110111_10001111_11110010;
assign in[613] = 496'b11111111_11111111_11111111_11111111_11111111_11111011_10001111_01000111_01001111_11001101_11111111_11011001_01000000_00010010_10101001_01110101_01010000_11111111_01001011_11001010_10111011_01001111_11000000_01101111_11110110_00110100_00110011_00001110_11101010_11111111_01001010_11111001_11111111_11111100_11111111_11111111_11110110_01001100_11111111_11111111_11111111_11111111_11111111_10111010_00101110_11111111_11111111_11111111_11111111_11111111_10010100_10110001_11111111_11111111_11111111_11111111_11111100_01010101_11100000_11111111_10110100_00100100;
assign in[614] = 496'b10111001_01101100_11111111_11111111_11111111_11111111_10100000_00111001_11111111_11111111_11111111_11111111_11111111_00100100_10110000_11111111_11111111_11111111_11111111_11101010_01101010_11110000_11111111_11111111_11110100_11111111_11010100_01000101_11111111_11111111_11111111_11111111_11111111_00000000_00000111_11111111_11111111_11101011_10100010_11111111_00100111_10100000_11111111_11110100_00110111_01011101_11111111_01001001_01001101_01001100_01110101_01111101_10010010_11111111_11110110_11101111_11101111_11101100_10001000_11111111_11111111_11111111;
assign in[615] = 496'b10010101_01111100_10100001_11111111_11111111_11111111_00010101_10000011_01000100_11111111_11111111_11111111_11111111_11111111_10011110_01101111_11111111_11111111_11111111_11111111_11111111_10011110_01110000_11111111_11111111_11111111_11111111_11111111_10011110_00110001_11111111_11111111_11111111_11111111_11111111_10011110_00100101_11111111_11111111_11111111_11111111_11111111_10011110_00110001_11111111_11111111_11111111_11111111_11111111_10000101_10001110_11111111_11111111_11111111_11111111_00000101_01000100_10111010_11111111_11010011_01011110_11000110;
assign in[616] = 496'b11011001_01011010_11101100_11111111_11111111_11111111_00000011_00011110_11111111_11111111_11111111_10111100_00111010_01111101_01101101_01010010_00111000_10110011_11111111_10101101_01101101_11010010_11011011_00010001_01111101_11111111_10000110_00111011_11111111_11111111_10010100_00111100_11111111_01001001_00001011_11111111_11111010_01011111_10111101_11111101_01010100_11001100_11111111_10010011_01011110_11111011_10001100_01101000_11111111_11111111_01011110_00000111_11111111_00101011_00101100_11111111_11111111_00111010_11010000_11111111_11111111_11111111;
assign in[617] = 496'b11111111_10010001_01100111_11111001_11111111_10000011_11111111_10000010_00001010_11111111_11111111_11111111_11111111_11110100_01010111_11010111_11101010_11000100_11110100_11100010_00011010_01111101_01100111_01100000_01111011_10001001_00000001_01110011_10001110_11100010_11011000_01111001_11111111_10111010_01100111_11111110_11111111_00100010_00011110_11111111_00011000_00011110_11111111_11000001_01101010_11011111_11010110_01110001_10110100_11110100_01001000_10100100_11111111_10100111_00100011_11111110_00101100_01011000_11111110_11111111_10110001_11000110;
assign in[618] = 496'b00000100_01100010_01111110_01111110_01110110_01011111_01101100_00001101_11100010_10100011_01111110_00111101_01001011_11101000_11111111_11111111_11101000_10110000_01111001_10000001_11111111_11111111_11111111_11111111_11111111_00100001_01110100_00101010_10001101_11001001_11111111_11111111_11111100_10010001_01010101_01111110_01101110_11111011_11111111_11111111_11010100_01100100_01101001_10100101_11111111_11111111_11011101_01110010_01000000_11101001_11100101_10001101_00111101_10101110_01111110_01011010_01010101_01111110_01110001_00000000_10001111_11001010;
assign in[619] = 496'b01011001_10100100_10100100_10010110_00010011_11110111_01011011_11111110_11111111_11111111_11111111_11111111_11111111_00001001_10101111_11111111_11111111_11111111_11111111_11111111_11110011_00001110_00001001_11010011_11111111_11111111_11111111_11111111_11101110_10010111_01000110_11100100_11111111_11111111_11111111_11111111_11111111_00110110_10111000_11111111_11111111_11111111_11111111_10100010_01101011_11010001_01000000_00101101_00010110_00000001_01100010_10010111_11111111_10101111_10101111_10000111_01000100_11010011_11111111_11111111_11111111_11111111;
assign in[620] = 496'b11111111_00011110_11111111_11100000_00111110_11111111_11111111_01000111_11111010_11111111_01000011_11111111_11111111_11111111_00101000_11010110_00100010_00101010_11111111_11111111_11111111_00010100_01110001_00000010_11111110_11111111_11101101_00011000_00110010_01101000_11011010_11111111_11010101_01001110_10110111_11111100_10000001_01001011_11111101_00000101_10000110_11111111_11111111_11110111_00100000_11111011_00100000_11100111_00010011_10110110_00101100_10111101_11111111_01100110_01111010_01000111_10011110_11100001_11111111_11111111_11111111_11111111;
assign in[621] = 496'b11111111_11111111_11100110_10010111_00000000_11001101_11111111_00001110_00101010_10101111_10010010_11111100_00101010_00111111_01011011_11110111_11111111_11000111_11111111_10101110_01111000_00111100_01000001_00111011_01011010_11111111_00011010_00010101_11111111_11111111_11111111_11111111_11111111_00010011_10010011_11111111_11111111_11111111_11111111_11111000_01111001_10010011_11111111_11111111_11111111_11111111_11111001_01110101_10010011_11111111_11111111_11111111_11111111_11111111_00000010_00100101_11011010_01000000_00001111_01110011_01111011_01100000;
assign in[622] = 496'b11111111_11111111_11111111_11111111_11111111_00100111_01101111_01000011_01100101_01000010_11110100_01100010_00100110_11110100_11111111_00011010_01101000_00010010_01000010_11110111_11111111_10110100_10001110_11001000_00110111_00011001_11100110_00000010_00110101_11111101_11011001_01100010_00110100_01010101_10001111_11111101_11111111_10011010_01011110_11111111_11111111_11111111_11111111_11111110_00111011_00110000_11111111_11111111_11111111_11111111_11011000_01111101_10110001_11111111_11111111_11111111_11111111_10000111_01110011_11111111_11111111_00010111;
assign in[623] = 496'b01000101_00001110_01001110_11100000_11111111_10001110_11111111_11111111_10100100_10100001_11111111_10010100_00000110_11111111_11111111_11001100_10000011_11111111_11111110_00010110_10111101_11111111_10100101_10110000_11111111_11111111_11111101_00111000_00010101_00100100_11110100_11111111_11111111_11111111_11110110_00000001_01110101_11110001_11111111_11111111_11111111_11111111_00000111_10100111_00011000_11101010_11111111_11111111_10010110_00000110_11111111_11100001_00001000_11111111_00000011_00111010_01100001_00001001_00111011_11111111_11010010_10110110;
assign in[624] = 496'b11101100_00000001_01001100_01011010_00110110_11100101_01100100_00101000_11010101_11111111_11110011_11111111_10001100_01000010_11111111_11111111_11111111_11111111_11111111_00010111_00100010_11111111_11111111_11111111_11111111_11111111_11100010_01100100_10000111_10100111_10001100_10010110_11111111_11001110_01011010_01010000_01000111_01110011_01111110_10111101_01100000_10101101_11111111_11111111_11110100_11010101_01001101_11000010_11111111_11111111_11111111_11111111_11111111_01001000_11000000_11111111_11110110_11010101_11111111_00110100_00110010_11001010;
assign in[625] = 496'b11111111_11111111_01110001_01001001_11111111_11111111_11111111_11111111_01111100_00101001_11111111_11111111_11111111_11111111_11010010_01111100_10101101_11111111_11111111_11111111_11111111_01000100_01011101_11111010_11111111_11111111_11111111_10011100_01111010_10100110_11111111_11111111_11111111_11110001_01010011_01101010_11111111_11111111_11111111_11111110_00100111_01111000_11001001_11111111_11111111_11110101_11110100_01110110_01111001_00100110_00100101_01001101_01011110_11111111_11000001_10000010_10000001_10000010_11000000_11111111_11111111_11111111;
assign in[626] = 496'b11101110_11111111_11111111_11111111_11111111_01011010_11001010_11111111_11111111_11111111_11111111_11111111_00000011_00000000_11111111_11111001_11111000_11111011_11111111_10100100_01100011_00110110_01001100_00011010_01010101_11111111_11000101_01111101_00111011_11111000_11111111_10100111_11111111_11000101_01111101_10110001_11111011_11111111_10101010_11111111_10101110_01111101_00101001_11000001_11111111_00011001_11111111_10010110_01111101_00101110_11001111_00110001_00100101_11111111_11111100_10100001_10000001_10000001_10111000_11111111_11111111_11111111;
assign in[627] = 496'b11100010_10011110_00001100_00111110_01111000_10010101_01011111_01000110_10100111_11000100_11011111_00110001_01111101_00000111_11110110_11111111_11111111_11111111_01111101_00100110_11101111_11111111_11111111_11111111_11101001_01111101_11000111_11111111_11111111_11111111_11111111_11010001_01111101_11000111_11111111_11111111_11111111_11010000_00111100_01111101_10111111_11111111_11111111_11001100_01000101_00000101_01110011_00111010_10101000_00101111_01010110_01111101_01111101_11001100_00101100_01101001_01111101_01111101_01101001_11101010_11011111_11011111;
assign in[628] = 496'b11111111_11111111_11111011_10101010_10000010_00000010_10111101_11010001_01001101_10010110_10110010_10001110_10011001_00110110_01110111_01110001_00010100_10011101_11111111_11111111_00011101_10110011_11010001_10100101_10001110_11111111_11100011_00110100_11111100_11111111_11111111_11111111_11111111_00000000_10101010_11111111_11111111_11111111_11111111_11111001_01011001_11010100_11111111_11111111_11111111_11111111_11101000_01011110_11111101_11111111_11111111_11111011_11111111_11110010_01101111_11010000_11000101_01010010_11001111_01010100_01111001_10010111;
assign in[629] = 496'b10111110_10000010_10000011_10000011_10101001_01011101_01101100_00100101_10010010_00110001_01111100_01100000_01101111_10101111_11111111_11111111_11111110_00011111_01111011_10011111_11111111_11111111_11111111_11111111_01001101_01111011_11010000_11111111_11111111_11111111_11111100_01010011_01111100_11010000_11111111_11111111_11111111_10101011_01111101_01111011_10001100_11111111_11111111_11111101_01001100_01110001_00111100_01000000_11011110_11001111_00111100_01111100_10010101_11110111_00110111_01101100_01101101_01101100_00001111_11111111_11111111_11111111;
assign in[630] = 496'b11111111_11111111_11111111_11111111_11111111_00111111_01111100_01111101_01111100_00101010_11010111_01110010_01010100_00000001_00010110_01111101_01111101_01011001_00011011_11111111_11111111_00011010_01100011_10011010_01111100_10001111_11111111_10101110_01101110_00011011_10111000_01111101_01111100_01111101_01110111_00000110_11111111_10101110_01111100_10111101_10010011_11001100_11111111_11111111_00111001_01001010_11111111_11111111_11111111_11111111_11011101_01111100_00010001_11111111_11111111_11111111_11111111_00011111_01111100_11001000_00110100_01110111;
assign in[631] = 496'b11111111_11110110_10100111_10100111_11110110_11111111_10001101_01100110_01100110_01100110_01010001_11110100_01000001_01111010_00000100_11110110_10110011_01111100_10010100_01111110_10000100_11111111_11111111_10111000_01111101_01100010_01001111_11111011_11111111_11111111_10000101_01100110_01111101_10000100_11111111_11111111_11101111_01101011_00110101_01111100_10010100_11111111_11111111_10010000_01111100_10111000_01101101_10000100_11111111_11100010_01111100_01000100_11111111_10101011_01110000_00110110_01101011_01111010_00101000_10010110_10010110_11010001;
assign in[632] = 496'b11111111_11101111_10100001_11111111_11111111_11100001_00110011_01110001_01111101_10110100_11111111_11011110_01011110_00001101_11100101_01111101_01010010_11111111_00010110_00010010_11110010_00110001_01011100_01011101_11111111_00100110_00101100_01010111_00010001_10000111_01010000_11111111_11101100_10110010_11011110_11111111_01001001_00000111_11111111_11111111_11111111_11111111_11111000_01110011_11000011_11111111_11111111_11111111_11111111_11000010_01110001_11101011_11111111_11111111_11111111_11111111_00100100_00010101_11111111_11011001_01110110_11000011;
assign in[633] = 496'b11111111_11001111_01101100_00110001_11111111_11111111_11111001_01101000_00100100_11010001_11111111_11111111_11111111_11010111_01101001_10000101_11111010_11111111_11111111_11100011_00001110_11110001_10101111_00110010_11011001_11110111_00000010_11001011_11111111_11111111_10111100_00110100_10101010_00000111_11111111_11111111_11111111_11101010_00111001_00110001_10110001_11110011_10011111_00100101_01011010_10011011_10100000_00001001_10000010_01111011_00101101_10101111_11111111_11111001_00010100_11010111_11000011_11111111_11111111_11110100_11111111_11111111;
assign in[634] = 496'b11111111_11111111_00000010_00110000_11111111_11111111_11111111_11000111_01110111_11010111_11111111_11111111_11111111_11111100_01001001_00000001_11111111_11111111_11111111_11111111_11000000_01010010_11110011_11111111_11111111_11111111_11101011_01101010_11000000_11111111_11111111_11111111_11111111_00111001_00000110_11111111_11111111_11111111_11111111_10100100_00110001_11111110_11111111_11111111_11101101_11110101_10001010_01000111_00010110_00001110_00111011_01110010_10000100_11001100_10010100_10011001_10100101_11010000_11111100_11111111_11111111_11111111;
assign in[635] = 496'b11111111_01001110_10100110_11111111_11111111_11111111_11111010_01101101_11101010_11111111_11111111_11111111_11111111_10111011_00110111_11111111_11111111_11111100_11111111_11110011_00010000_01000010_00011101_01001011_01000111_10110011_10101000_01110011_10010111_11101010_11000110_00110010_11111111_11110001_01011110_11110100_11111111_00000011_10111100_11111111_10111101_00011011_11111111_11111111_01000110_11110001_11000000_00101011_11010101_11111111_00010100_10001101_11111111_10100101_01010010_11111001_11111111_00010110_11110010_11111111_11111111_11111111;
assign in[636] = 496'b01010100_01001110_00101011_01100011_10010110_11111111_11111111_11111111_11101011_01101010_11010110_11111111_11111111_11111111_11111001_01000000_10010110_11111111_11111111_11111111_11111111_00001110_00100011_11111111_11111111_11111111_11111111_00000000_00110001_11111111_11111111_11111111_11111111_00010101_00111000_11110010_11111111_11111111_11111111_10100100_01001110_11110010_11111111_11111111_11111111_11111001_01100011_11011101_11111111_11111111_11011101_00000111_01101010_01110001_00011100_00111000_01110001_01111000_00110001_10110010_10111001_11110010;
assign in[637] = 496'b11011100_00010010_00011001_10001101_01000110_11111111_00001100_11100100_11111111_11111111_11111010_11111111_11111100_00011000_11111010_11111111_11111111_11111111_11111111_11110010_01010011_11000010_11111111_11111111_11111111_11111111_11111111_11000101_01010101_01010000_00110010_11010100_11111111_11111111_11111111_11101101_11010111_10101110_10011110_11111111_11111111_11111111_11111111_11111101_11010100_11110110_11111111_11111000_10111100_00001101_00010100_11010001_11111111_00011001_01011010_00101000_00100011_11010100_11111111_11111111_11111111_11111111;
assign in[638] = 496'b00000101_11100001_11111111_11111111_11111111_11111111_00101010_11101010_11111111_11111111_11111111_11111111_11111111_00110001_11110010_11111111_11111111_11111111_11111111_11111110_01001100_11111001_10100100_00110011_00110100_11111111_11111011_01011100_01000110_00000000_11101010_10100001_11111111_11110100_01111110_10010111_11111111_11111111_00001010_11111111_11110100_01110100_11101001_11111111_11001111_01000000_11111111_11010001_01111110_10011110_00010110_01001001_11010111_11111111_11111111_10100001_10000001_10110001_11110101_11111111_11111111_11111111;
assign in[639] = 496'b11011000_01001000_01100111_01011000_01011010_11000010_01101000_00010000_11110010_11100110_01001111_11100110_01010111_10001000_11111111_11111111_10101101_01011111_00000110_01000010_11111110_11111111_11111111_00101001_01010011_01000101_11000110_11111111_11101011_10011101_01100101_10011000_01011110_11001100_11111111_10100100_00100111_01111101_11101111_01010101_11101000_11111111_10100100_01111101_00010111_11111111_00110001_11001100_11111111_00100100_01111101_10010101_11111111_10010001_00010111_00001011_01111001_00010101_11110110_10000001_11000101_11111111;
assign in[640] = 496'b01111100_01110101_00111010_11001100_11111111_00101011_11111111_10111100_01110101_10011100_11111111_10010011_00110001_11111111_11100001_11011101_11111111_11111111_11111000_01101010_10001011_11000000_10111000_11111111_11111111_11111111_11001011_01111100_01111110_00011100_11111111_11111111_11111111_11011000_01111110_10001010_11111111_11111111_11111111_11111111_10110101_01111110_11100010_11111111_11111111_11111111_11111111_11011000_01111110_11001100_11111111_11101111_10001011_11111111_11110111_01001110_01110000_01000101_01110111_11100101_10011110_10100001;
assign in[641] = 496'b01010000_10111011_11111111_11111111_10011110_10000101_00000000_11111111_11111111_11111111_11110001_11111111_00010100_10111101_11111111_11111111_11111111_11111111_11111111_11001001_00001010_11111111_11111111_11111111_11111111_11111111_11111111_00100010_01000000_00101110_11111111_11111111_11111111_11111111_10001000_00111000_10111100_11011011_11110001_11111111_11011000_01000001_11110101_00011001_01100000_00000011_11111111_00010000_10100111_10011110_01111101_01100110_11100100_11111111_10000011_01111110_01000001_00111110_10110011_11111111_11111111_11111111;
assign in[642] = 496'b01111100_11100101_11111111_11111111_11111111_00111011_01110111_11101100_11111100_11000001_11010010_11100111_01110100_01111001_00011000_01101110_01111101_01110001_10001011_01111101_01101011_01111101_01000100_00000110_01111011_10001010_01101001_10010001_11010101_11111111_00100011_01111101_11111111_11111111_11111100_10101010_00111011_01111101_01001110_11111100_10011011_00000011_01110110_01111101_01110000_10111110_10001001_00011010_00100010_01111001_01100000_11011101_11111111_00010111_01110111_01111101_01010110_11011101_11111111_10000101_11101100_11111111;
assign in[643] = 496'b11111111_11110011_00101100_11111111_11111111_11111111_11111111_11101110_01001100_11111111_11111111_11111111_11111111_11111111_10111001_00011111_11111111_11111111_11111111_11111111_11111111_00000001_00010000_11111111_11111111_11111111_11111111_11111111_00110111_10111010_11111111_11111111_11111111_11111111_11111111_01000000_11101111_11111111_11111111_11111111_11111111_11111111_01011110_11111111_11111111_11111111_11111111_11111111_11000100_01011000_11111111_11111111_11111111_11111111_11111111_10100011_10000011_11111111_11111111_10010110_11000100_11111111;
assign in[644] = 496'b00011011_00011100_11010001_11100000_10011000_11110101_00101110_11111110_11111111_11111111_11011011_11111111_11111111_00110000_11111100_11111111_11111111_11111111_11111111_11111111_11010011_00010111_10101100_11010001_11111111_11111111_11111111_10110100_01011001_01010001_01111100_11011001_11111111_11010000_01001001_11101001_11111110_11100000_11111011_11111111_00101100_10110111_11111111_11111111_11111111_11111111_11111111_01010011_11111000_11111111_11011110_10000010_11111111_11111111_10000011_00101100_00100001_01110111_00111100_10001101_10111010_11101101;
assign in[645] = 496'b11111111_11111111_11111111_11111111_11111111_11101111_00010110_01010001_00011001_10110101_11111111_11111111_00011000_10011100_11111111_10001101_01011101_11111111_11111111_00011010_10001001_00111001_10100101_01010100_11111111_11111111_11110001_11000111_11110011_11111111_00110110_11111111_11111111_11111111_11111111_11111111_10111110_00000000_11111111_11111111_11111111_11111111_11111111_00010000_11010100_11111111_11111111_11111111_11111111_11111111_00101110_11111111_11111111_11111111_11111111_11111111_10110100_10001000_11111111_11111111_00100001_11101010;
assign in[646] = 496'b11000111_00110110_01110101_01111101_01111101_01000110_01110000_00101010_10010110_10101001_10001101_01010110_01010110_11001010_11111111_11111111_11111111_11111111_00111100_11101110_11111111_11111111_11111111_11111111_11110110_11001010_11111111_11111111_11111111_11111111_11111111_10011010_11111010_11111111_11111111_11111111_11111111_10111111_01110100_11111111_11111111_11011011_10011100_10100010_01011111_01101101_11101001_11111111_00001100_01111110_01111101_01110001_10111110_01101011_01001110_01101000_01111100_00101010_11101011_10000001_11000010_11111111;
assign in[647] = 496'b11111111_11111111_11111111_11111111_11111111_10111000_01100100_01110001_01011010_01101100_01111100_11010101_01101101_11000100_11111001_10001011_01110100_01111100_11100011_01011110_01101011_01011101_01111110_01111110_00010010_11111111_11111000_11011110_11001011_10010001_01111101_11000110_11111111_11111111_11111111_11111010_01011010_00111111_11111111_11111111_11111111_11111111_00010011_01110111_11001010_11111111_11111111_11111111_11001100_01111011_00000010_11111111_11111111_11111111_11110001_01011001_01000001_11111001_11111111_01000101_11101001_11111111;
assign in[648] = 496'b11111111_11111111_11000100_10011101_11111111_11111111_11111111_10111010_01111101_01110111_11111111_11111111_11111111_11111111_01000010_01111110_00101000_11111111_11111111_11111111_11111111_01001101_01111110_10111110_11111111_11111111_11111111_11111111_00011000_01011100_11111011_11111111_11111111_11111111_11010101_01101101_11011110_11111111_11111111_11111111_11111111_00101010_00010010_11111111_11111111_11111111_11111111_10101100_01101100_11011001_11111111_11111111_11111111_11111111_01011001_00011000_11111111_11111111_11111111_11101011_11111111_11111111;
assign in[649] = 496'b01011010_01100111_01000011_10010111_11111111_01110010_00111000_10001001_10010100_01011000_10111010_00001100_11101100_11111111_11111111_11111111_11110101_11111010_01000010_10100100_11110100_11110111_11110011_11110011_10101111_01100001_01111101_01111001_01100100_01111101_01111101_01111101_11110111_11100010_10010100_10010100_10010100_10010100_01010101_11111111_11111111_11101110_11101001_11101001_11000111_00111101_11001110_00110111_01101111_01111101_01111101_01111101_01111101_11111111_11001001_10011101_10011101_10011101_10011101_11111111_11111111_11111111;
assign in[650] = 496'b11111010_00110001_01111100_01011111_01100110_11111111_10010000_01110001_10110100_11111100_01000111_11111111_11111111_01000101_00010101_11111111_11111111_00110001_11111111_11111111_01011000_10000001_11111111_11011001_01110010_11111111_11111111_00010101_01010000_10110110_01100010_10000010_11111111_11111111_11100011_01111110_01111101_00110010_11111111_10111001_00101111_01011100_01000110_01111000_01100101_11110101_00111111_01111101_00110110_11010001_01111000_01111001_11001110_00000101_01111101_01100001_01111100_01101001_10110000_10010011_10100001_11110110;
assign in[651] = 496'b01111101_01001011_11111111_11111111_11111111_11110110_01111101_00100010_11111111_11111111_11111111_11111111_10100101_01111101_10111001_11111111_11111111_11111111_10100101_01101001_01111101_10100101_11001101_11000011_11000011_00000100_01111101_01111101_01111101_01111101_01111101_01111101_10101111_01111101_01001011_10101111_00011000_00011000_01111101_01000001_01110011_11110110_11111111_11001110_00100011_01110011_01110011_10101111_11111111_11111111_10000110_01110011_00100010_11010111_11111111_11111111_11111111_00001110_00110110_11111111_11111111_11111111;
assign in[652] = 496'b11111111_10000101_01111100_01111010_01111101_11111111_11111111_11001111_11010011_11011011_00010101_11111111_11111111_11111111_11111111_11011011_00111100_01111101_11111111_11111111_11101010_00010110_01101111_01100001_10111111_11111111_00001010_01101111_01110001_10001011_11110101_11111111_00111000_01111101_00110010_11010110_11111111_11111111_11111111_01111011_10001001_11111101_11111111_11111111_11111111_11111111_01110111_10001110_10110010_11010010_11111111_11101011_11111100_01110001_01111101_01111101_01111100_01011100_01110010_11001010_10111111_10001001;
assign in[653] = 496'b11111111_11010111_01110100_00001110_11111111_11111111_11111101_00110110_01010011_11111001_11111111_11111111_11111111_10001011_01111000_11001010_11111111_11111111_11111111_11100000_01110010_00010000_11100100_11000011_11111101_11111111_00010010_01111110_01010000_01111011_01110100_00011110_11011001_01110011_00101011_10110110_11101011_00110110_00101001_10110101_01111110_11001011_11111111_10011111_01111001_11000000_10111011_01111110_00110000_00110111_01110101_00000011_11111111_10110011_01100110_01010101_00100110_11001101_11111111_11111111_11111111_11111111;
assign in[654] = 496'b11111111_11100101_01111110_10100101_11111111_11111111_11111111_10000010_01111100_11100001_11111111_11111111_11111111_11111111_00111001_01100001_11111111_11111111_11111111_11111111_11111111_01011100_00010010_11111111_11111111_11111111_11111111_11101001_01111101_10010001_11110010_11111111_11111111_11111111_10100111_01111110_10011011_11111111_11111111_11111111_11111111_00010110_01111110_00100110_11111111_11111111_11111111_11111111_00011011_01111110_10111011_11111111_11111111_11111111_11111111_10001010_01110011_11110110_11111111_11011110_10010011_11111111;
assign in[655] = 496'b10101011_11111111_11111111_11111111_11111111_00110101_11100000_11111111_11111111_11111111_11111111_10110001_01110001_00110101_11100110_11111111_11111111_11111111_01111100_01111101_01110010_10110001_11111111_11111111_11111111_00011011_01001101_11111000_11111111_11111111_11111111_10111100_00001001_00001000_11111111_11111111_11111111_11111111_11111111_10000101_01101111_00011101_00001000_00001010_00100000_00011001_11110010_10010110_00101100_00110011_01001000_00111101_01001001_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111;
assign in[656] = 496'b10101010_01010000_01111001_01110010_01111100_10000110_01110010_01010101_10100101_11101001_00011010_10100000_01111011_00100111_11110101_11111111_11111111_10110000_00100010_01110100_11100101_11111111_11111111_11111111_11110101_01111001_00110011_10100110_00100001_01101011_01101010_00110001_01111110_01111101_01111110_01000110_10000001_10000010_00111110_01111101_01011101_10100101_11111111_11111111_11111111_00011100_01110001_01001011_11110101_11111111_11111111_10100110_01111100_10111110_01110001_01011111_00100010_00110001_01110101_10010001_10000010_10000001;
assign in[657] = 496'b10111100_10010110_11100110_11111111_11111111_00011001_01000000_00011001_01100101_10011000_11111111_11111111_01110001_11100010_11111111_10101000_01110100_11001111_11111111_00110011_10010011_11010011_01011100_01000100_10100001_11111111_11100001_00101110_01001100_10111101_10000110_10100001_11111111_11111111_11111111_11111111_11111111_00111011_11001101_11111111_11111111_11111111_11111111_10101110_01010000_11110110_11111111_11111111_11111111_11010111_01011100_11000001_11111111_11111111_11111111_10010100_01100011_11010001_11111111_01001101_11101011_11111111;
assign in[658] = 496'b01010100_01101110_01111010_00111011_11101000_11001011_01111101_11001001_11000000_01001100_10001000_11111111_11001011_01110011_11111101_11111111_11111101_11111111_11111111_11001011_01110110_11110001_11111111_11111111_11111111_11111111_11001011_01111011_01010011_00111110_11100010_11111111_11111111_10111110_01111101_01110111_01101010_01000001_11111111_11111111_10010000_01111101_10100101_00011011_01111000_11111111_11111111_10011110_01111101_10111000_01110001_01110001_11111111_11111111_10110111_01111101_01110001_01110100_10111011_10111010_10000001_10100110;
assign in[659] = 496'b11111111_11111100_11000110_01111100_01001100_11111111_11111111_11110110_00010111_01111100_00111100_11111111_11111111_11111111_11010000_01111100_01111100_11000110_11111111_11111111_11111111_00100010_01111100_00110000_11111110_11111111_11111111_11100111_01110110_01111101_10110010_11111111_11111111_11111111_10000010_01111101_01010000_11111111_11111111_11111111_10101011_01101000_01111101_10101000_11111111_11111111_11111111_01000000_01111100_01011011_11111111_11111111_11111111_11111111_01010100_01111100_11000000_11111111_11111111_10100111_11111111_11111111;
assign in[660] = 496'b11010001_00100100_01010011_01011000_10011110_00010111_01111011_01111101_01111101_01111101_01111001_00111001_01111101_01010100_10010010_11011010_01110011_01111101_01111101_10001010_00010001_01001011_11010001_01111101_01111101_01111101_10001100_11101101_01010010_01011111_01111101_01111000_01111010_01100101_10111001_10011101_01111101_01111101_01011101_00000001_01111101_01111101_00101101_01111101_01111101_10011010_11111000_00100100_01111101_01111101_01111101_01001101_11101011_11111111_11010110_01110010_01111101_01111101_10101000_01110101_00001101_11001010;
assign in[661] = 496'b11010111_10000111_10000011_10111101_11110111_00011010_01110111_01111100_01111011_01111011_01010100_11100011_01111010_01010000_10011100_10100001_01010101_01111101_11110111_01011100_01111011_00110010_10110110_01101000_01101011_11111111_10111110_01010011_01111011_01111011_01111011_01000100_11111111_11111111_11111111_11010011_01111100_01101101_11011010_11111111_11111111_11111111_10001111_01111011_00000101_11111111_11111111_11111111_11111111_01010000_01110011_11101000_11111111_11111110_11111010_10110001_01110111_00010100_11111111_01111011_01010000_11111111;
assign in[662] = 496'b11101000_00110000_01111001_01001101_11000110_11111101_01000011_10010000_11101011_11000001_01000101_11111111_11100110_00101110_11111111_11111111_11111111_10100000_11111111_11110001_01011011_11110001_11111111_11111111_11111111_11111111_11111111_00001100_00101100_11111100_11111111_11111111_11111111_11111111_11111001_01010001_01011000_01010111_10111011_11111111_11111111_11111111_11111100_11110110_00001001_11000011_11111111_11111111_11111111_11111111_11100011_00101001_11111100_11100000_10001111_00011011_01001110_01001011_10111001_00000101_11000010_11111110;
assign in[663] = 496'b11111011_01100001_10100111_11111111_11111111_11111111_10111101_01110111_11110011_11111111_11111111_11111111_11001111_00010110_00111100_11111111_11111111_11111111_10101000_01100000_01111110_10000001_11111110_11000100_00101010_11111111_11011000_01111110_01000101_01011000_01011110_01111110_11111111_10101110_01111010_00011111_11000101_10010011_01011011_11111111_10000111_00100001_11111111_10110011_01101101_11001110_11111111_01000101_10101111_11111111_10001000_10101110_11111111_11010000_01110001_11110001_11111111_11111111_11111111_11111111_11111111_11111111;
assign in[664] = 496'b01111000_01000001_00000110_11111111_11111111_00110100_11100010_11111111_11111111_11111111_11111111_01101100_00100111_11000101_11110100_11111111_11111111_11111111_11001000_01000000_01110100_01101101_00001001_11111010_11111111_11111111_11111111_11101111_10111011_01111101_10110110_11111111_11111111_11111111_11111111_10100111_01100111_11110010_11111111_11111111_11111111_11100100_01011111_00000110_11111111_11111111_11111111_11111111_00001000_01111101_00001001_00001001_10100000_11111111_11111111_10110101_00010110_00010110_00010110_11111111_11111111_11111111;
assign in[665] = 496'b11111111_11111111_00110010_00101110_11111111_11111111_11111111_10011011_01101011_11100100_11111111_11111111_11111111_11101001_01100100_10011000_11111111_11111111_11111111_11111111_00101100_01000011_11110011_11110001_11100011_11111111_00001010_01111101_01001001_01011000_01110110_01010010_00111111_01011011_10110110_11110110_11111111_11110001_01010001_10010010_11110101_11111111_11111111_11111010_10101000_01101101_00001000_10101011_00010000_01000001_01100111_01010110_10110010_10110111_10000001_10000001_10110001_11011100_11111111_11111111_11111111_11111111;
assign in[666] = 496'b11111111_00001000_10000010_11111111_11111111_11111111_11111111_01010101_10110111_11111111_11111111_11111111_11111111_11100011_01110111_11011001_11111111_11111111_11111111_11111111_11000111_01100010_11111101_11111111_11111111_11111111_11111111_10011010_00110100_11111111_11111111_11111111_11111111_11111111_10000101_00001011_11111111_11111111_11111111_11111111_11111111_00100010_00001011_11111111_11110110_11111111_11111111_11111111_00010101_01110100_01101011_01101111_00100100_11111111_11111111_11110100_10100011_10000010_10101011_11111111_11111111_11111111;
assign in[667] = 496'b11101010_11110011_11111111_11001100_00010001_01010001_01111100_01101111_01011010_01110110_01111101_11111111_00000001_01000001_00110101_01111110_01010111_11010000_11111111_11111111_11010110_01100100_01000000_11101101_11111111_11111111_11110011_01001011_01000100_11110010_11111111_11111111_11111111_10010101_01110000_11011011_11111111_11111111_11111111_11111111_01011110_00001000_11111111_11111111_10110100_00110011_11111111_01100111_10011010_11111111_11101011_00111110_01101100_11111111_01100110_00101010_00011111_01100110_01101000_01111101_01110011_10010000;
assign in[668] = 496'b11111111_11111111_11111111_11111111_11111111_10010000_01000100_01100010_00100111_11001000_11111111_00100001_01011001_10110010_10101011_00111011_01111000_10110101_01101010_11101011_11001111_01100101_11000011_00101000_00110001_01111010_01011000_01111101_01001011_11101110_10011011_01101110_10100110_00000011_10010110_11101111_11111111_10011011_01111101_11111111_11111111_11111111_11111111_11111111_10011010_01100110_11111111_11111111_11111111_11111111_11111111_00010011_00110100_11111111_11111111_11111111_11111111_11100001_01110111_11111111_11111111_00010000;
assign in[669] = 496'b01111101_01110110_01000101_11101101_11111111_01111101_00011011_10000100_01110011_01000010_11111111_11110000_01001010_01110100_10110100_10101001_10100011_11111111_11111111_10110100_01111101_01110100_10100001_11010011_11110101_11111111_11111111_10000011_01111101_01111101_01111010_01001011_11111111_11111110_00100000_01111101_01101110_00001110_00001110_11111111_10101110_01111101_01011011_11001010_11111111_11111111_11111111_11101000_01111101_01100101_00000010_11010010_11000100_11111111_11111011_00010001_01101010_01111101_01111101_11111111_11110011_11001110;
assign in[670] = 496'b10000010_10101011_11100000_11111111_11111111_01111101_01111101_01111101_01111101_00011000_11111111_01000111_10000111_00011010_01111101_01111101_01111101_10000100_11000111_11111111_10010000_01111101_01000001_01111000_01110001_00101111_00101010_01111001_01101111_11110001_01001100_01111101_01111101_01111101_01111101_00001101_11111111_00010110_01111101_10010000_00001100_11001000_11111110_11111111_01101111_01111101_11111111_11111111_11111111_11111111_11011010_01111000_01111101_11111111_11111111_11111111_11011001_00110010_01111101_10011010_01111011_01111101;
assign in[671] = 496'b01100100_11111001_11111111_11111111_11111111_01011010_01111110_11110000_11111111_11111111_11111111_11111111_01111011_01111111_11110000_11111111_11111111_11111111_11111111_01111011_01111110_11110000_11111111_11111111_11111111_11111111_01111011_01010101_11111110_11111111_11111111_11111111_11011101_01111101_00011000_11111111_11111111_11111111_11111111_11000010_01111110_00101010_00001100_00001100_00100100_01001101_11100011_01111100_01111101_00111111_00111011_00010010_10000111_11111111_11100011_11101110_11111111_11111111_11111111_11111111_11111111_11111111;
assign in[672] = 496'b01011100_01110001_01111011_01101110_00110101_00111101_00011010_00101001_00110010_01111100_01111101_11111111_11111111_11111111_11110111_00110001_01111011_01001110_11111111_11111111_10100101_01100101_01111011_01011011_11010010_11111111_10100100_01110110_01111101_00100110_11100000_11111111_10111001_01110110_01111011_10001000_11110110_11111111_11111111_10010010_01111101_00010001_11111111_11111111_11111111_11111111_10110000_01111100_01001111_10011101_10100010_00011001_01010101_11111000_00100111_01101110_01111100_01111011_01111011_11100101_10110111_10110011;
assign in[673] = 496'b00111101_00111110_01000001_01101110_00011101_00011101_11111111_11111111_11111111_10110101_01100000_00111101_01111100_10111110_11111111_11111111_11110111_10110001_10001100_01110111_01101100_11001000_11111111_11111111_11111111_11111111_10001010_01110111_01101110_01001000_10101011_11111111_11111111_00000001_01110111_01111100_01100100_10100100_11111111_11001011_01111010_01101001_10011100_11110110_11111111_11111111_10110001_01111010_01101000_00101101_11000000_11110001_11010100_11111111_10100101_01011010_01111100_01111011_01111011_11110100_10110111_10000010;
assign in[674] = 496'b01010011_01100011_01111101_01011001_10010100_11111010_11111111_11111001_10010111_01111000_01111100_11101110_11111111_11111111_11111111_11111111_00011101_01111101_11101110_11111111_11111111_11111111_11111111_10011000_01111101_10110011_11111111_11111111_11111111_11111111_10011000_01111101_01100110_11010110_11111111_11111111_11111111_00000010_01111101_01110011_01110110_00100101_10000110_01011110_01111010_01111101_10111000_01011011_01111101_01111101_01111101_01111101_10001100_11111111_00001011_01111101_01111101_01101000_10011000_10010000_10111010_11101010;
assign in[675] = 496'b01101111_01111111_01111111_01111111_01101111_01111111_01111111_00000000_11000000_00000000_01101111_01111111_01010000_11100000_11111111_11111111_11111111_11010001_01111111_11010001_11111111_11111111_11111111_11111111_11111111_00110000_11111111_11111111_11111111_11111111_11111111_11010000_10100000_11111111_11111111_11111111_11111111_11111111_10010000_10010001_11111111_11111111_11110000_11111111_11000000_01111111_01010000_00000000_00000000_01100000_01100000_01101111_01100000_01111111_01111111_01111111_01011111_01111111_00100000_11000000_11111111_11111111;
assign in[676] = 496'b11111111_11111111_11111111_11111111_11111111_01101000_11100100_10001101_00010101_00010101_00000100_10011110_01111101_01111011_01111001_00111001_00011110_01011110_10111000_01111101_01111101_01101111_01000011_00100010_10001001_10111000_01101101_11011101_10011011_00100010_00111101_00111101_10111000_01111101_11001001_11111111_11111111_11111111_11111111_10111000_01111101_10001101_11111111_10111011_11101101_11111111_10111000_01111101_00011000_11011110_01101011_00001110_11111111_11111011_01001001_01111010_01000000_01111101_10001010_01101111_01111101_01001110;
assign in[677] = 496'b11110011_10000100_01101010_00111110_10111100_11111110_01000101_01111110_01011000_01000110_01111000_11011000_01001010_01101010_00001100_11111001_11111110_01011111_01010001_01111110_00011010_11111111_11111111_11111111_01011001_01111110_00100111_11111000_11111111_11111111_11111000_01110011_01111110_11010110_11111111_11111111_11111111_11001011_01111110_01111100_10100100_11111111_00001000_10011111_01101011_01100001_00100101_01000110_11111111_00011011_01111110_00101111_11010011_10111000_01111011_00000001_01100101_00100011_11111111_01010111_01000011_11100010;
assign in[678] = 496'b01010011_01001101_00100001_10110001_11111011_11111011_01010001_01111101_00101011_01011000_00111001_11111111_11111111_10010110_01111101_10101101_11111010_10111010_11111111_11111111_11111001_00110011_01101110_00000000_10101100_11111111_11111111_11111111_11111001_00110000_01111100_01111101_11111111_11111111_11111111_11111111_11111111_10101011_01111101_11111111_11111111_11111111_11111111_11111111_11100010_01111101_10101011_10011101_00100001_00101000_11010101_11000111_01011010_01111011_01111001_01011011_00001001_11100101_11101001_11111111_11111111_11111111;
assign in[679] = 496'b11111100_11111111_11111111_11111111_11111111_01111111_11101100_11111111_11111111_11111111_11111111_00110111_01111111_11101100_11111111_11111100_10100010_10111101_00110111_01111110_11100111_10001100_01011110_01111110_01111110_10000010_01111110_01000100_01111110_00111010_10101101_01111110_11010100_01111010_01111110_00000001_11111001_00000011_01111110_11111111_01101110_00111101_11110111_10101001_01111110_01010000_11111111_10000100_01110111_01011110_01111110_00111101_11011110_11111111_11011011_01010100_00111100_10101100_11110111_11111111_11111111_11111111;
assign in[680] = 496'b01101100_11110000_11111111_11111111_11111111_00100001_01100001_11111111_11111111_11111111_11111111_11111011_01011010_01011001_11111111_11111111_11111111_11111111_10111000_01111110_10001100_11111111_11111111_11111111_11001010_00011010_01111101_11110010_11111111_11111111_11110111_01101101_00011010_01111101_11101110_11111111_11111111_11101111_01111101_11000011_01110001_01010111_00110010_00100101_00101000_01111110_11111111_11110101_10000001_00011011_00011011_01101010_01111101_11111111_11111111_11111111_11111111_11111111_00011010_11111111_11111111_11111111;
assign in[681] = 496'b10010110_11111111_11111111_11111111_11111111_10110000_00010000_11111111_11111111_11111111_11111111_11111111_00101011_11000100_11111111_11111111_11111111_11110001_11010100_01010110_10100010_00000000_00110010_01111010_01111101_00100011_00111011_00101001_00101001_00001010_11000001_01001000_01000101_11111110_11111111_11111111_11111111_10000111_00011010_00111100_11111111_11111111_11111111_11110100_01010101_11101110_00001000_11111111_11111111_11111111_10010110_00010001_11111111_11100110_11111111_11111111_11111111_00010011_11000001_11111111_11111111_00011010;
assign in[682] = 496'b11000101_10001111_10101111_11100101_11111111_10001000_01111001_01111101_01111100_01110100_01010000_11111111_01100001_01001110_11011111_11011111_11000011_10011100_11111111_01001101_01110111_10011000_11101011_11111100_11111111_11111111_11011100_01110011_01111110_01100000_01101010_10110010_11111111_11111111_11100101_10000010_01010011_01111100_00001100_11110010_11011111_11001011_10011101_00111101_01111100_00000110_01101001_01111100_01111100_01111101_01111100_01100000_11101101_10001111_10001111_10100100_11010001_10000001_10111011_11111111_11111111_11111111;
assign in[683] = 496'b11110101_11010100_00010110_00110011_00001001_10000110_01011111_01111110_01111101_01111101_01111101_00111110_01111101_01111000_01100000_00100100_00101111_01110111_01111101_00000101_11011011_11111111_11111111_11111111_00001101_00000101_11111100_11111111_11111111_11111111_11111111_00001101_10111101_11111111_11111111_11111111_11111111_11001000_01110010_00110001_11110111_11111111_11110100_00000001_01100100_01111101_01111101_01011101_00100100_01100010_01111101_01111101_00110100_01000100_01111101_01111101_01111110_01111101_00111110_00110001_00011110_10010001;
assign in[684] = 496'b10011010_01111110_10111101_11111000_11111111_11000011_01101011_01111111_01111110_10010001_11111111_11111111_11111111_10101101_01111110_10001011_11110101_11111111_11111111_11111111_11001001_01111111_11011101_11111111_11111111_11111111_11111111_10110000_01111011_11100001_11111111_11111111_11111111_11111111_10000100_01011101_11111111_10110111_10110000_11111111_11111111_10000100_01011101_00010100_01110010_10001101_11111111_11111111_10000100_01111100_01100011_11100100_11111111_11111111_11111111_10000111_01111110_10101110_11111111_11110100_10110011_11111000;
assign in[685] = 496'b10011111_01111001_10110010_11111111_11111111_11111111_10001011_01001011_11110001_11111111_11111111_11111111_11111010_10001101_00110111_11111111_11111111_11111111_11111111_11001000_01111101_00010000_11111111_11111111_11111111_11111111_10001010_01111000_10110110_11111111_10111100_11100111_11111111_00000110_01100001_11111111_11111111_01010100_00110100_11111111_10111001_01101111_11011100_11111111_00000111_01111110_11111111_11011110_01100111_01110101_00000001_01011011_01110111_11111111_11111111_11110000_10001000_01000010_01111101_11111111_11111111_11111111;
assign in[686] = 496'b11111111_11111111_11111111_11111111_11111111_10001001_01011011_01001100_10001000_11111111_11111111_00100010_00011000_11110100_11111000_00001010_10000110_11111111_01100101_11111011_11111111_11010101_00000001_01000111_11111001_01010000_00010110_00001000_01100110_10000100_00110010_11001101_11111111_10110111_10011111_11100100_11111111_00101111_11000000_11111111_11111111_11111111_11111111_11111111_00010101_11000000_11111111_11111111_11111111_11111111_11111111_00110010_11000111_11111111_11111111_11111111_11111111_11110110_01001110_11111111_11111111_10111000;
assign in[687] = 496'b11111111_11000001_10001000_11100111_11111111_00111110_00101101_01111101_01111101_01111100_01010010_11111110_01110001_01111101_00010000_11100111_11000110_01000000_11101010_01110110_01111101_10001110_11111011_11110010_00100001_11001100_01111101_01110100_01111101_01101001_01101110_01100110_11100000_01111001_10011000_11011011_11000011_10100110_11110011_11111111_01101011_00101100_11111111_11111111_11111111_11111111_11111111_00000110_01110111_11000101_10010010_11000000_11111111_11111111_11100000_01110101_01011110_01110111_00000011_10001011_01111101_01111101;
assign in[688] = 496'b11111111_11111111_11111111_11111111_11111111_11111111_11000100_01100100_01001111_00100101_11101000_11111111_11111111_10101001_01000011_11100001_01100110_11000011_11111111_11111111_11110110_01011100_01110001_10011000_11111111_11111111_11110101_00111000_00000001_00000000_00110011_11110011_11111111_00000101_00010010_11111111_11111111_00001001_10100000_11111111_01100111_11011101_10100011_00100110_01010100_10101110_11111111_01010111_11111111_11111000_10101101_11010111_11111111_11101100_00110010_11111111_11111111_11111111_11111111_11111111_11111111_11111111;
assign in[689] = 496'b11101010_10011010_10000010_10111000_11111111_10101001_01110001_00111001_00010111_01101010_10100101_10100101_01000001_11001000_11111111_10000011_00100111_00110001_10100101_01010011_00101011_00110010_01100110_01010111_00011000_11111111_11010000_10101010_11001110_11010011_01110101_11010011_11111111_11111111_11111111_11111110_00111011_00110100_11111101_11111111_11111111_11111111_00010100_01100000_11100111_11111111_11111111_11111110_00010011_01101101_11010101_11111111_11111111_11110101_00100001_01010111_11010110_11111111_11111111_11101000_11111111_11111111;
assign in[690] = 496'b11000111_10101010_10011000_11111011_11111111_10001111_01011111_10100101_10001011_00100011_11011110_11111111_11111111_00001011_00111110_11101000_01000101_10110110_11111111_11111111_11111100_00001011_01110010_00110001_11111111_11111111_11111111_11111111_00000010_00111111_01010101_11101110_11111111_11111111_10010001_10011010_11111111_10010111_00100010_11111111_10001000_00011110_00111111_10001101_01100010_00011111_11110111_01100011_11010001_11010000_10101111_10110111_11101011_10100111_01000001_11111111_11111111_11111111_11111111_11111111_11111111_11111111;
assign in[691] = 496'b11111111_11001101_10101010_11101000_11111111_11111111_11111111_10100011_00111110_00011010_00000101_11111111_11111111_11111111_11110010_01001101_00011011_01100111_11111111_11111111_11111111_11011000_01100011_00011101_11111010_11111111_11100110_00111010_00011010_11110000_00100100_10111010_11111111_00111010_00010010_11011001_10011001_10010110_01000101_11000001_01001110_11111100_11111111_00010010_00100001_11011010_00100011_10011000_11111111_11111111_11111111_11111111_11111111_01000010_11110010_11111111_11111111_11111111_11111111_11111111_11111111_11111111;
assign in[692] = 496'b11111111_11111111_11111111_11111111_11111111_01010110_01110010_00110000_00010101_11110011_11111111_00101001_11101000_10010101_01111101_01111101_00100000_11111111_11001101_11111111_10110000_01111101_01010010_01100111_11011111_01110111_01110110_01111011_01100111_11101010_01111101_00010111_10011110_01010101_01001100_10101110_11111100_01011110_01001000_11111111_11111111_11111111_11111111_11111111_01001001_00110110_11111111_11111111_11111111_11111111_11001000_01111101_10000101_11111111_11111111_11111111_11111111_00010101_01111101_11111111_11100001_01110110;
assign in[693] = 496'b01000000_11111111_11111111_11111111_11111111_10100000_01101111_11111111_11111111_11111111_11111111_11111111_11110000_01111111_11110000_11111111_11111111_11111111_11111111_11111111_01100000_10010001_11111111_11111111_11111111_11111111_11111111_01000000_00101111_10010001_01100000_00000000_11111111_11111111_01000000_01111111_01111111_01010000_01000000_11111111_11111111_00110000_01010000_11110000_00011111_00010000_11111111_11111111_11100000_01111111_01010000_01111111_11010000_11111111_11111111_11111111_00010000_01111111_00000000_11111111_11111111_11111111;
assign in[694] = 496'b11111111_11111111_11111111_11111111_11111111_10010000_11110101_11101100_10110110_00001001_10010110_11111100_00110010_01101100_01110000_00000011_00001010_00001101_11101001_01101001_10011100_00110111_01010001_11011001_11111111_10001011_00011110_11111111_11111111_10011111_01010011_10000110_00011010_10101101_11111111_11111111_11111111_11010101_10010000_00100111_11101100_11111111_11111111_11111111_11111111_11111111_00110011_11000000_11111111_11111111_11111111_11111111_11111111_00011010_00011000_11111111_11111111_11111111_11111111_11000101_11111111_11111111;
assign in[695] = 496'b11111111_11111111_11111111_11111111_11111111_00010001_01001110_01011101_01110000_00111100_11010101_01000010_10101111_11101101_11111111_11110110_10010110_01101000_11011001_11111011_11011001_10001100_00101000_00001110_00001111_01010011_01010011_00110001_10011001_10111010_11111111_10000100_11111111_11111111_11111111_11111111_11111111_11111111_00100101_11111111_11111111_11111111_11111111_11111111_11001111_01010100_11111111_11111111_11111111_11111111_11100010_01011101_10101001_11111111_11100001_11111111_11101000_01010010_10000001_10110000_01010001_00000010;
assign in[696] = 496'b10111101_00101011_01110101_01111101_00111111_00000111_01111000_00111100_10000110_10100001_01011101_10100100_01110011_10101110_11111111_11111111_11111111_11001101_01000000_10000101_11111111_11111111_11111111_11111111_11110111_01110001_11011101_11111111_11111111_11111111_11111111_10101011_01110001_11101110_11111111_11111111_11111111_11111101_01000010_01100010_11111111_11111111_11111111_11111111_00000101_01101101_01111001_11100000_11111111_11111101_00001000_01111000_10101000_01111101_10000100_00001100_01011000_01111001_10011101_01000111_00101000_11011101;
assign in[697] = 496'b01101111_01111111_11000000_11111111_11111111_00100000_11111111_10010000_01111111_10010000_11111111_10110000_00000000_11111111_11111111_00010000_01111111_11111111_11000000_00010000_11111111_11111111_00000000_01111111_11111111_11110000_01111111_11010000_11111111_00000000_01111111_11111111_11111111_00010000_10110000_11111111_00000000_01111111_11111111_11111111_11010000_01101111_11110000_01100000_01100000_11111111_11111111_11111111_01000000_01011111_01111111_10110000_11111111_11111111_11111111_10110000_01111111_01000000_11111111_11111111_10010000_01011111;
assign in[698] = 496'b00001101_00000010_01101001_10000011_11111111_00111010_11111111_11111111_11101010_01100011_11101100_10100101_01001011_11111111_11111111_11111111_01100110_11100100_11100100_01110101_10011110_11111111_10101001_01101100_11110010_11111111_10110000_01101111_00100111_01101001_10111110_11111111_11111101_10101000_01001101_01011011_01010101_11010001_11111111_11110111_00011010_11110010_11110010_00001111_01100101_10110100_11001000_01010101_11111111_11111111_11111111_11011100_01101001_11001000_01111000_00111010_00011010_10001011_00011010_10011010_10000010_10000001;
assign in[699] = 496'b01001001_01111100_01111011_01010100_00001011_01100111_01001011_01001100_01011100_01111011_01111011_01010001_11100100_11111111_11111111_11101111_01000111_01111011_11010101_11111111_11111111_11111111_11111111_11010000_01111011_10010101_11111111_11111111_11111111_11111111_11110101_01010110_01011100_11101111_11111111_11111111_11111111_10001110_01111011_01111011_00100010_11010000_00110110_01110001_01111011_01111011_01000111_01111011_01111011_01111100_01111011_01111010_01101111_11110000_00101000_01111011_01111100_00000100_10111001_11001001_10001100_11111000;
assign in[700] = 496'b11010101_10001111_10100010_11111110_11111111_00110101_00100011_10110010_00000010_01000010_11100100_00010001_10001111_11111111_11111111_11111111_10001110_00001100_01001001_11110111_11111111_11111111_11111111_11111011_01010100_00011110_11111111_11111111_11111111_11111111_11111111_00010001_00101111_11111111_11111111_11111111_11111111_11111111_00010111_01000111_11011001_11111111_11111111_11111111_11111111_01000011_11001111_00101011_11110101_11111111_11111111_11101100_01001110_11111111_11000011_00000001_11111111_11111111_10000101_11111111_11101000_10110001;
assign in[701] = 496'b11111111_11100000_01111100_10001010_11111111_11111111_11111111_00011100_01100010_11101101_11111111_11111111_11111111_11010010_01110100_10011000_11111111_11111111_11111111_11111000_01001000_01010101_11111101_11111111_11111111_11111111_00000100_01111011_11000111_11111111_11111111_11111111_11010010_01111101_10000010_11111111_11111111_11111111_11111111_01000000_01101111_11000100_11011111_11101100_11011111_11111001_00100000_01111101_01111101_01111010_01110101_01111010_01101110_11111111_11110011_10111110_10111110_10111101_10111110_11111111_11111111_11111111;
assign in[702] = 496'b01110000_11101000_11111111_11111111_11111111_00101101_01111101_11011101_11111111_11111111_11111111_11111111_10010110_01111101_00011101_00001110_00001110_11000001_11111111_10000110_01111101_01000000_10101011_00011110_01101001_11111111_00101101_01111101_00111101_11111111_11110111_01011110_11111111_00101101_01111101_01110010_11110110_11111111_00111011_11111111_10000001_01111101_01111101_10100100_00100111_01111001_11111111_01010010_01111101_01111101_01111101_01111101_00110100_11111111_11101101_11000001_10000001_10000001_10100010_11111111_11111111_11111111;
assign in[703] = 496'b10111101_10010011_11111111_11111111_11111111_11111111_00011000_11000000_11111111_11111111_11111111_11111111_11111101_01010001_11111001_11111111_11111111_11111111_10011000_10001010_01010011_10011000_10001110_11111100_11111111_11000001_00000111_00010111_10110000_10111110_11111111_11111111_11111111_00010010_00100010_10010000_10101000_10111110_11110001_11111111_10110000_11001001_11001001_10100011_10000010_00100000_11111111_11111111_11111111_11111111_11111111_11111111_11011000_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111;
assign in[704] = 496'b00001110_00011100_11111111_11111111_11111111_11111111_00100101_10010111_11111111_11111111_11111111_11111111_11111111_01101011_11001010_11111111_11111111_11111111_11111111_11100111_01111011_10001001_11000000_11111100_11111111_11111111_11011011_01110001_10011111_00111001_01010000_00010110_11111111_11000001_01000100_11111111_11111111_10110100_01111110_11111111_00001110_10000011_11111111_11110111_01011010_00101011_11111111_00110101_11001011_11111111_10010100_01011110_11110100_11111111_11111101_11111111_11111111_01011101_11000100_11111111_11111111_11111111;
assign in[705] = 496'b01001101_01110011_01101110_01100000_01111001_01110111_01000111_11001000_11101010_11111010_10111110_00011010_01111101_11001100_11111111_11111111_11110011_10001010_11001000_01111101_01111100_00111100_10010110_00110010_01111000_11111111_11001010_01111100_01111101_01111101_01111101_00100111_00011011_01101000_01111100_01001111_10000010_01010111_01110000_01111010_00000010_11101110_11110010_11111111_11001101_01111101_11000000_11110000_00000001_10010010_10001010_00111001_00101100_01011100_01101011_01000110_00101111_00101111_10010010_11110000_11111111_11111111;
assign in[706] = 496'b11111111_10101011_01111000_11100111_11111111_11111111_11111110_01000101_10001000_11111111_11111111_11111111_11111111_10101100_01100100_11111010_11111111_11111111_11111111_11111111_00111010_00001010_11111111_11111111_11111111_11111111_11110011_01111001_01000011_01011010_10101001_11111111_11111111_00010011_01100111_10011100_10110110_01110001_11100101_11111111_01110001_11001001_11111111_11111110_01100010_11011010_11111111_01110001_11111000_11101110_00011110_00011110_11111111_11111111_00101101_01110000_00001101_10110111_11111111_11111111_11111111_11111111;
assign in[707] = 496'b11111111_01100111_11111111_11111111_11111111_11111111_11111100_01100110_11111111_11111111_11111111_11111111_11111111_11111100_01100111_11111111_11111111_11111111_11111111_11111111_11101011_01010010_11111111_11111111_11111111_11111111_11111111_11010010_00100100_10101000_10110100_11111111_11111111_11111111_10110000_01111011_00000010_01000111_11101101_11111111_11111111_00100100_10000110_11111111_00101010_11101001_11111111_11110010_01110001_11101111_11110000_01011110_11110011_11111111_11110110_10100010_10111101_01010010_10110100_11111111_11111111_11111111;
assign in[708] = 496'b11111111_10100110_10001001_00111010_10100001_11111111_11111111_00000000_11111111_00001110_10011100_11111111_11111111_11111111_10101111_10001010_01010010_11111010_11111111_11111111_11111111_11101111_01111000_10111111_11111111_11111111_11111111_11111111_10001010_01100100_11001101_11111111_11111111_11111111_11000110_11001100_00011010_10111000_11111111_11111111_11111001_10001110_11111111_00100001_11110001_11111111_11111111_00001011_11100101_10111110_00000001_11111111_11111111_10111110_10010101_10111001_00110001_11110011_11111111_00001001_11110110_11111111;
assign in[709] = 496'b11111111_11111111_11011101_11010110_11111111_11111111_11111001_00100001_01100001_01000010_01011010_11111111_11111111_10010100_01000000_11110110_11111111_11111100_11111111_11111111_10100000_01101111_01000100_00011010_11000110_11111111_11111111_11111111_11110010_10111100_01110101_10101011_11111111_11111111_11111111_11111111_10001001_01000100_11111111_10101101_10000101_01001010_01000001_01010100_11101111_11111111_00110010_10010101_10111111_00010000_11100011_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111;
assign in[710] = 496'b11010001_00111100_01111101_01111101_01000010_11100010_01100100_01001111_10111001_10010011_01111101_11111111_10011001_01111101_11011010_00000001_01111000_01000010_11111111_10010101_01111101_01011110_01011010_10010100_11111100_11111111_10001101_01111101_01111101_01011000_11000110_11111111_11101111_01101011_00010010_00001011_01100011_01111011_00010010_10000011_01000101_11111101_11111111_11101101_01000011_01110100_01100101_00010011_11111111_11101000_10011111_01110110_00111001_10110010_01011000_00001000_01100010_01110011_00100010_01111110_00111101_11101111;
assign in[711] = 496'b11111111_10000101_01010101_11111010_11111111_11111111_11101101_01011010_10101011_11111111_11111111_11111111_11111111_00000111_00111110_11111101_11111111_11111111_11111111_11000000_01101010_10100011_10011000_10110000_11111011_11110001_01011111_01111010_00100110_00100010_01001000_00011011_00100100_01111110_01000101_11111111_11111111_11001101_01010110_10100010_00100111_00000101_11111111_11111111_00100000_00001111_11111111_01001001_00001010_10001011_00110101_00101001_11111001_11111111_11011010_10001001_10000111_11001000_11111111_11111111_11111111_11111111;
assign in[712] = 496'b11111111_11110000_10010001_01000000_00110000_11111111_11010001_01100000_01010000_00010000_00100000_11111111_11000000_01101111_10100000_11111111_11111111_11111111_11010001_01101111_10010000_11111111_11111111_11111111_11111111_01010000_00101111_11111111_11111111_11111111_11111111_11110000_01101111_11100000_11111111_11111111_11111111_11110000_01010000_00000000_11111111_11111111_11000000_11000000_01100000_01010000_00100000_11000000_10110000_01101111_01111111_00010000_11111111_01111111_01111111_01101111_00100000_11000000_11111111_11111111_11111111_11111111;
assign in[713] = 496'b11111111_11111111_11101010_10001011_10001011_00000001_11101100_11001011_01100100_00100110_01100100_00000010_00011100_01101101_01110001_00000101_11101010_01101011_11111111_11111111_01010001_01011111_01011111_01100000_10101000_11111111_10111101_01100011_11101001_11110101_11101111_11111111_11111111_00010011_00011010_11111111_11111111_11111111_11111111_11111111_01000001_10001110_11111111_11111111_11111111_11111111_11111111_00110010_10101010_11111111_11111111_11111111_11111111_11111111_00001010_00011110_11111111_11011110_00101110_01101111_00100001_01101111;
assign in[714] = 496'b11111111_11101110_01011100_11111111_11111111_11111111_11111111_10001011_00110110_11111111_11111111_11111111_11111111_11110000_01010001_11000111_11111111_11111111_11111111_11111111_10001000_01010011_11111111_11111111_11111111_11111111_11111000_01101011_10110110_11000111_10011000_11011001_11111111_00001011_01001111_01000110_00101110_10001000_01010111_11111010_01011111_01100101_10110010_11111111_11000010_01101100_11100011_10001011_00101000_00011011_00110011_01101100_10110111_11111111_11111111_11100110_10000001_10010101_11100011_11111111_11111111_11111111;
assign in[715] = 496'b11111111_11111111_11111111_11111111_11111111_11101010_10001110_10000001_10000001_10100000_11010010_00010011_01111100_01000100_00111100_01111110_01100101_01111010_01010101_10101111_11110010_00011000_01011110_11110000_00010001_11001001_11111110_10000110_01000010_11010011_11001111_01100100_01110010_01100100_00001001_11101010_11101010_01100010_01000001_11011110_11101100_11111111_11111011_00111111_01011111_11011000_11111111_11111111_11111111_00000101_01111110_11000101_11111111_11111111_11111111_10111100_01110011_10011011_11111111_01010110_10010001_11111111;
assign in[716] = 496'b11111111_11111111_11110001_01000101_01111101_11111111_11111111_11010101_01001101_01111101_01100101_11111111_11111111_11100100_01011011_01111101_01111101_10101010_11111111_11111101_01000111_01111101_01111011_10011000_11111111_11111111_00001001_01111101_01101011_10110001_11111111_11111111_11011111_01101011_01111101_10010000_11111111_11111111_11111111_11000000_01111101_01010101_11111101_11111111_11111111_11111111_11110000_01101101_00110101_11111111_11111111_11111111_11111111_11111111_11001010_00110110_00010110_00010011_00010011_11111111_11001001_10001010;
assign in[717] = 496'b11111011_10111100_10110100_10110111_11110001_11100000_01100010_01111001_00110010_01011101_01111001_11111111_00100001_01010111_11010101_11111111_11111111_10101111_11111111_10011000_01111000_10001100_10111010_00100000_01100001_11101010_10001010_01111111_01111111_01111110_01010100_10101011_01100101_00110011_10111001_11100010_00100010_01110011_11011000_10000011_11111101_11111111_11111111_11111110_00110101_00101111_11111111_11111111_10110001_10010110_10100101_01101010_10001001_00110001_01011011_01010101_01010101_01001001_11001001_11111111_11111111_11111111;
assign in[718] = 496'b11111111_11111111_11111111_11111111_11111111_00001101_00101100_00111110_00111001_11111000_11111111_00001100_11001011_11111111_11111111_01010001_10000111_11111111_00011010_11110001_11111111_11110010_01001001_00111101_11111111_11001000_00111001_10111110_00111000_10101011_01000000_11111111_11111111_11011001_10010110_11011111_10111110_00001000_11111111_11111111_11111111_11111111_11111111_00001001_11000100_11111111_11111111_11111111_11111111_11111111_00101100_11111011_11111111_11111111_11111111_11111111_11001111_10000011_11111111_11111111_00010000_11101001;
assign in[719] = 496'b11010101_01101100_01110111_01111101_11001111_11101111_01011101_00110000_11100100_00000011_11010101_11111111_00011010_01000110_11111011_11111111_11111111_11111111_11110000_01111001_10101000_11111111_11111010_11100110_11111111_11101100_01100011_10011011_11010100_01011011_01000111_11111111_11111111_10100001_01111011_01111011_01111101_00101011_11111111_11111111_11111111_11000110_10101101_01110101_10001111_11111111_11111111_11111111_11110101_10101111_01111001_10010000_11111111_11010011_10001111_01101100_01111101_01011010_10100110_10010101_11000111_11111110;
assign in[720] = 496'b11111111_10100000_00000000_10100000_11111111_11110000_01010000_01101111_00110000_01111111_10110000_11111111_00010000_01010000_11110000_11111111_01010000_00000000_11111111_01101111_11000000_11111111_11111111_01010000_00000000_11111111_01010000_00101111_10110000_01010000_01111111_11100000_11111111_11010001_00110000_01000000_01101111_01100000_11111111_11111111_11111111_11111111_11010000_01111111_11000000_11111111_11111111_11111111_11111111_01010000_00100000_11111111_11111111_11111111_11110000_00101111_01100000_11110000_11111111_01000000_11110000_11111111;
assign in[721] = 496'b00100001_00111001_10100101_11001010_00000110_10001000_00011000_11111111_11111111_11111111_11111111_11111111_01000110_11011000_11111111_11111111_11111111_11111111_11111111_00011110_11010011_11111111_11111111_11111111_11111111_11111111_10111110_00110011_11111100_11111111_11111111_11111111_11111111_11111111_10010001_00101000_11000110_11110010_11111111_11111111_11111010_10110101_00100100_01111110_01010011_11111001_11001010_01011110_00010010_11001000_11111001_11111111_11111111_10001110_00110110_00101010_00111010_00000101_11111111_10000001_10100100_11110101;
assign in[722] = 496'b11001001_00101111_00101111_10000111_11110001_11111111_00011100_01010111_10011101_10010100_10000010_11111111_11111111_10110101_01111101_10001010_11111100_11111111_11111111_11111111_11111111_10011101_01110010_10000001_11111111_11111111_11111111_11111111_11111111_11001110_01100011_00010010_11111111_11111111_11111111_11111111_11111111_11100110_01100100_11111111_11111111_11111111_10110000_10001001_10001001_01101001_10101011_00010100_01010011_01001110_00011011_00011011_00000011_00101111_10010101_11010100_11111010_11111111_11111111_11111111_11111111_11111111;
assign in[723] = 496'b11111111_11111111_11111111_11111111_11111111_10100111_11100001_10010000_00010101_10100001_11111111_10101010_01100100_01100111_00011011_10010100_01111110_11001010_11111111_11001110_01111100_01000100_00000111_00001000_11111100_11111111_11010110_01111001_11010111_11111111_11111111_11111111_11111111_11110101_01011100_00010011_11111110_11111111_11111111_11111111_11111111_10111100_01111010_00010000_11111110_11111111_11111111_11111111_11111111_10100001_01101010_10100011_11111111_11111111_11111111_11111111_11111111_10100101_01110100_11111111_11111111_11111111;
assign in[724] = 496'b11111111_11111111_11010111_01000010_01100101_11111111_11111111_10100110_01010101_11000010_00100101_01011011_11101110_11010111_01100100_11011101_11010101_01011111_01000001_00101101_01010011_10110111_10111001_01010000_10110110_11101000_00111000_01111101_01110000_01001011_11001100_11111111_11111111_10000101_00110111_11100000_11111111_11111111_11111111_11111111_10000101_00000110_11111111_11111111_11111111_11111111_11111111_10000101_00010101_11111111_11111111_11111111_11110010_11111111_10110100_01101000_11000111_11011100_10001010_10001001_01100010_01111110;
assign in[725] = 496'b11111111_11111111_11111111_11111100_11000100_01111101_10110000_11111111_10111000_01100001_01101111_11111100_00101011_01100100_00110110_01111010_00101110_11100101_11111111_10101011_01111101_01111101_01111101_01110101_01100010_11011001_01111101_01011100_10101111_10100001_10001101_10110110_10000011_01110110_11100100_11111111_11111111_11111111_11111111_01100111_10001000_11111111_11111111_11111111_11111111_11111111_01110001_10011100_11111111_11111111_11111111_11111111_11111111_00011100_00110111_11111111_11101101_10101111_11000001_01001000_01110010_00101011;
assign in[726] = 496'b10111001_01000011_01011111_00100100_01000011_10101010_01111100_00101110_11111001_11111111_11110010_11111101_01001111_01100101_11111001_11111111_11000100_01100101_11111010_01100000_01101011_10001001_01000001_01000100_10101010_11111111_11100000_01110111_01111100_01111101_01001101_11011100_10011111_01100101_00011011_11011100_11010011_01000110_01000100_01101100_10000010_11111111_11111111_11111111_11000000_01101001_00010110_11111111_11101101_10001011_10001110_01101001_10010001_00101111_01000110_01101111_00111101_00011011_11000111_11110011_11111111_11111111;
assign in[727] = 496'b11111111_11111111_11011101_01010001_10011100_11111111_11111111_11110101_01000010_00011101_11111111_11111111_11111111_11110111_00111101_00101100_11110101_11111111_11111111_11111111_00101100_01011011_11100001_11111111_11111111_11111111_10000001_01111001_10111111_11111111_11111111_11111111_11100101_01100100_00000000_11111111_11111111_11111111_11111111_00011010_01110100_11110100_11111111_11111111_11111111_11111111_10000010_01110100_00011110_10100001_00000110_10001110_00011010_11111111_11000101_10000010_10000001_10000010_10000010_11111111_11111111_11111111;
assign in[728] = 496'b01011111_11111111_11111111_11111111_11111111_11010101_01100001_10101010_11111111_10110000_00100011_11111111_11111111_10010110_01100100_01000100_01101001_10010000_11111111_11110011_00001100_01101100_01011000_01110011_01010101_11110110_00111111_01010110_11100000_11111111_11101011_11111001_00100110_01100110_11101000_11111111_11110111_00000100_11101011_01110001_00001110_11111111_11111111_11111111_10111011_11101110_01111100_11011011_11111111_11111111_11111111_11111111_11111111_00011010_01010001_10101110_11101010_11100111_11110000_01000111_01111101_01111110;
assign in[729] = 496'b11111111_11111111_11010011_11010000_11110100_11111111_11011100_01001001_00100100_00100001_01011001_11111111_11111111_00001011_10000110_11111111_11111111_10111001_11111111_11111111_10100000_01001011_10001010_10100110_11011101_11111111_11111111_11111110_11001100_00011110_01111011_01000111_11111111_11111111_11111111_11111111_11110011_01011101_11100011_11111111_11101111_11001001_00010101_00101000_10011000_11111111_01010011_01011000_00101110_10110000_11100111_11111110_11111111_11111010_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111;
assign in[730] = 496'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11101001_10100101_01001011_00011011_00111011_10101000_00010001_10010000_00010000_00011011_11111011_11111011_10011001_11111011_11100011_00110011_11100011_11111111_11111111_11011010_10011110_01010001_11010001_11111111_11111111_10011011_00001100_11011001_11111000_11111111_11111111_10001001_10010001_11111111_11111111_11111111_11111111_10111010_00000010_11111111_11111111_11111111_11111111_11111111_11111000_11110010_11111111_11111111_11111111;
assign in[731] = 496'b11111111_11111111_11111111_11111111_11111111_10000100_10001011_11001000_11101101_11110011_11111111_01111101_01111101_01111110_01111101_01111101_01100101_00101111_11101100_11101100_11101100_10001011_10001011_01010100_01111101_11111111_11111111_11111111_11101010_00001111_01101100_01001010_11111111_11111111_11101010_01010111_01100011_00000000_11111001_11111111_11100111_01001111_00001001_11011100_11111111_11110110_11111111_01001011_01100000_11111111_10111111_00010001_01011001_11111111_01011011_01110110_01101001_01101000_01010111_11000101_11000101_11100000;
assign in[732] = 496'b00000011_01111101_01111100_01000010_11110101_01011001_01111100_01111101_01110001_01111101_10111010_00110000_01111101_01010011_11001000_11110111_11001000_11110001_01011110_01111100_11010000_11111111_11110110_11100101_11111111_10001111_01111101_01101111_01010011_01100011_01111110_11000110_11111111_11001110_00101010_01111101_01111100_01111101_10111010_11111111_11111110_00111110_01111101_01010001_11000101_11111000_11111111_11010110_01111101_01000011_11101101_11111111_11110001_11111111_11111110_00110111_01110110_01000000_00111100_11111010_00100011_01111101;
assign in[733] = 496'b11100001_01101111_10111010_11111111_11111111_11111111_11111111_01000001_10000001_11111111_11111111_11111111_11111111_11111111_01101010_10000010_11111111_11111111_11111111_11111111_11111111_01010110_00101000_11111111_11111111_11111111_11111111_11111111_01101010_01000111_11111111_11111111_11111111_11111111_11111111_01101011_00001010_11111111_11111111_11111111_11111111_11101001_01110010_11001010_11111111_11111111_11111111_11111111_11001010_01110010_11101001_11111111_11111111_11111111_11111111_10010111_01101011_11111111_11111111_00101000_00101101_11111111;
assign in[734] = 496'b11111111_11111111_11111111_11111111_11110000_01110010_10101010_11100000_00000101_01000101_01111010_11111111_10111101_01110011_01100011_01110011_10001111_10101001_11111111_11001001_01111100_01110100_01011010_00110110_01101110_11111111_01000010_00110000_11110111_11111111_11111111_11111111_11000110_01101111_11101110_11111111_11111111_11111111_11111111_10110011_01110000_11111100_11111111_11111111_11111111_11111111_11001110_01101011_11000111_11111111_11111111_11111111_11110101_11111111_01001111_00111010_11010001_10011100_00101011_01010010_01111110_01011000;
assign in[735] = 496'b11111111_00011000_01010110_11110111_11111111_11111111_11011100_01111011_11000101_11111111_11111111_11111111_11111111_00101001_00110101_11111101_11111111_11111111_11111111_11101000_01101010_00100001_00010100_00001111_11011111_11111111_00000001_01111101_01111101_00110001_00100000_01001101_11111111_01011001_01111101_00000010_11111110_11111111_01111000_11101011_01111101_01101100_11110001_11111111_10110101_01011101_11111111_10010101_01101011_00100000_01101001_01010001_11001101_11111111_11111011_10001011_10010010_11000101_11111001_11111111_11111111_11111111;
assign in[736] = 496'b11111111_11111111_11111111_11111111_11111111_11011010_00011001_01010001_01100100_01001111_10011100_10111101_01101010_10000100_10101011_01111110_00000100_01110010_01010011_10111011_11110011_01000000_10100011_10110110_01101010_01100010_10001111_01011001_10100111_11101011_01100101_10011110_10010001_00010011_11001100_11111111_00101100_00011111_11111111_11111111_11111111_11111111_10101001_01010010_11110111_11111111_11111111_11111111_11011010_01101001_11001110_11111111_11111111_11111111_11110100_01001111_10010000_11111111_11111111_01000000_11111110_11111111;
assign in[737] = 496'b11111111_11101101_00100100_01110010_01001000_11111111_11010000_01010011_00111101_10100100_10111110_11111111_11110001_01101011_00101101_11111010_11111111_11111111_11111111_10011000_01101010_11111010_11111111_11111111_11111111_11111111_10110100_01111011_00110111_10001101_10001101_11001110_11111111_11111111_00010100_01111000_01011001_01110011_01011110_11111111_00000101_01101001_10111010_11111111_11101100_11100101_11011101_01111101_10110110_11111111_11111111_11111111_11111111_11011000_01111010_00000011_11010110_10100111_10000011_01010110_01111101_00110100;
assign in[738] = 496'b11111111_11010001_01010100_11001000_11111111_11111111_11111111_10100111_01111101_11001101_11111111_11111111_11111111_11111111_00001101_01101100_11111111_11111111_11111111_11111111_11111111_00111100_00110101_11111111_11111111_11111111_11111111_11110001_01110010_10001101_11111111_11111111_11111111_11111111_11010011_01111110_10100010_11111111_11111111_11111111_11111111_11000100_01111110_10100010_11111111_11111111_11111111_11111111_10100010_01111110_10100100_11111111_11111111_11111111_11111111_10101011_01111110_10111111_11111111_11101001_01001111_11110100;
assign in[739] = 496'b11100111_10001100_00100010_10100100_11010111_10111010_00111000_10101010_11111111_11111111_11111111_11111010_00111000_11101110_11111111_11111111_11111111_11111111_11100111_01000010_11111111_11111111_11111111_11111111_11111111_11111111_10001011_00010101_11110110_11111111_11111111_11111111_11111111_11111111_10111100_00111000_11000000_11111111_11111111_11111111_11111111_11111111_11100101_00101110_11111011_11111011_11111111_11110001_10011000_01100000_01011110_00111000_01000011_10011111_00110011_00000111_10100101_11101111_11111111_11111111_11111111_11111111;
assign in[740] = 496'b11110110_10011101_00000111_00000111_10110001_10110011_00111100_10000101_10011100_10011100_00101111_01000000_00011111_11110101_11111111_11111111_11111111_11111101_00000101_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111010_11111111_11111111_11111111_11111111_11111111_11101011_00110101_11100110_11111111_11111111_11111111_11111111_00010011_10101000_01100000_00000001_11111111_11111011_10001001_01100001_11111111_11000100_01101101_11001110_00100001_01010100_00110110_01000011_10001110;
assign in[741] = 496'b11111111_11111111_11011010_10010110_10010110_11111111_11111011_00011100_01010010_00000101_10001000_11111111_11111111_00000100_00111101_11110011_11111111_11111111_11111111_11111111_01000101_10110100_11111111_11111110_11110111_11111111_11111111_10101000_01110011_01000010_01101010_00001100_11111111_11111111_11111111_11000111_00010000_01110011_11001111_00001001_00011001_00100001_01000011_01111101_10001110_11111111_10010101_10010101_11000000_10011001_10001100_11111100_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111;
assign in[742] = 496'b01011110_01110000_00111100_11110111_11111111_00011001_11111001_11101100_01010001_11001011_11111111_10000100_11100101_11111111_11111111_10110101_10001001_11111111_10100010_10000101_11111111_11111111_11011010_10000011_11111111_11111001_00110101_00010111_11111011_11000000_11000111_11111111_11111111_11111111_10001011_01001110_00011000_11110101_11111111_11111111_11111111_11110110_00101001_01110011_01010011_10001110_11111111_10101000_01011001_00101000_11111001_10111111_00100111_11111111_10111110_11010110_00100010_10010111_00001101_11111111_11000000_10100101;
assign in[743] = 496'b11111111_11111111_00101100_11011011_11111111_11111111_11111111_11101000_01100101_11111111_11111111_11111111_11111111_11111111_10101111_00111110_11111111_11111111_11111111_11111111_11111111_10100110_00010101_11111111_11111111_11111111_11111111_11111111_01000001_10110100_11111111_11111111_11111111_11111111_11111111_01110100_11100101_11111111_11111111_11111111_11111111_11111111_01011110_11111100_11111111_11111111_11111111_11111111_11111111_01011001_11111111_11111111_11111111_11111111_11111111_11111111_00111111_11111111_11111111_11111111_00000001_11111111;
assign in[744] = 496'b11111111_11111111_11111111_11111111_11111111_00000101_01101111_01111110_01010010_01011100_11000001_10011010_01100010_10110011_11010010_01011001_01101010_01110011_01010010_10011101_11000110_00100000_01000001_11100010_00000011_01010111_01110111_01000000_10010111_11111110_11110001_01011000_11101001_11010011_11111111_11111111_11100110_01001011_01001010_11111111_11111111_11111111_11010011_01011001_00111100_11101010_11111111_11111111_11100101_01011100_00010110_11110101_11111111_11111111_11100110_01011000_00100110_11111111_11111111_00111011_11110101_11111111;
assign in[745] = 496'b11111111_11111101_00001100_01001100_11101100_11111111_11111111_10010100_01010001_11110000_11111111_11111111_11111111_11100001_01011111_11010001_11111111_11111111_11111111_11111111_00101100_00011111_11111111_11111111_11111111_11111111_11000101_01101001_10011001_10011110_11011100_11111111_11101101_01010100_01110101_00000000_10111110_01101110_11101100_10001001_01001111_10101111_11111111_11010100_01101001_11110001_01010000_00000010_10011101_00010010_01110000_10111010_11111111_11001000_10000001_10000001_10111001_11110010_11111111_11111111_11111111_11111111;
assign in[746] = 496'b11111111_11110011_10110110_10011110_10011111_11110101_10001100_01101000_01111101_01111110_01111101_11111111_00101110_01101011_10000011_11010101_11111111_10101111_00110101_01011100_11010010_11111111_11111111_11111111_11010110_01011111_11110001_11111111_11111111_10101100_11101011_00000100_11010010_11111111_11111111_11111111_00110000_01001010_01111000_11111001_11111111_11101001_10000111_01111010_01111110_00111111_00100011_00100011_01100001_01111101_01111100_00011111_11111111_00101001_00101001_10000110_11100100_11100100_11111100_11111111_11111111_11111111;
assign in[747] = 496'b11110111_10010100_00011110_01101011_01111010_11011101_01010111_01100110_00100000_10010111_10110111_11111111_01000100_01010110_11101000_11111111_11111111_11111111_11101110_01110100_10100100_11111111_11110101_11111101_11111111_11111111_01000010_01100111_01010010_01111101_01011101_11111110_11010010_01001111_01100111_01001111_01000110_10010101_11111111_01010011_01001110_11011011_11111111_11111111_11111111_11111111_01111101_11001110_11111111_11111111_11110010_11111001_11111111_01000111_00101001_10011100_00010111_01110000_00111100_01100010_00100011_10110011;
assign in[748] = 496'b11111010_00010011_01111111_01100011_11100101_11111111_10000001_01111000_00111001_01111100_10010101_11111111_11101101_01111001_00010111_11111111_01101111_00010011_11111111_11010000_01111100_11000010_11111111_01101111_01011001_11111111_10101111_01110011_11110001_11011001_01110110_10010000_11111111_00010010_01000001_11111111_00110100_01111011_11100000_11111111_00010010_01110101_00000011_01111100_10011100_11111111_11111111_10001111_01111110_01111110_00010001_11111100_11111111_11111111_10110010_01111101_01001000_11111001_11111111_11001110_00101000_11110100;
assign in[749] = 496'b11111111_11111111_11111111_00011111_01111100_11111111_11111111_11111111_11010111_01110010_01111101_11111111_11111111_11111111_11110001_01101000_01110111_10111000_11111111_11111111_11111111_00001011_01111110_00000110_11111111_11111111_11111111_11010111_01111100_01001001_11111111_11111111_11111111_11111111_00100101_01111101_10011110_11111111_11111111_11111111_11001000_01110010_00111010_11111111_11111111_11111111_11111111_00101010_01111101_11010111_11111111_11111111_11111111_11110110_01111100_00110101_11111111_11111111_11111111_11100110_11111111_11111111;


    always @(posedge clk)
    begin
        if (read_input == 1'b1)
            out = in[addr];
        else
            out = 495'bZ;
    end

endmodule   
module get_label(input [9:0] addr, input read_input, output reg [3:0] out);
    
reg[3:0] label[0:749];

assign label[0] = 4'b1000;
assign label[1] = 4'b0110;
assign label[2] = 4'b0001;
assign label[3] = 4'b0100;
assign label[4] = 4'b0110;
assign label[5] = 4'b1000;
assign label[6] = 4'b1001;
assign label[7] = 4'b0100;
assign label[8] = 4'b0000;
assign label[9] = 4'b0101;
assign label[10] = 4'b0111;
assign label[11] = 4'b0100;
assign label[12] = 4'b0000;
assign label[13] = 4'b0101;
assign label[14] = 4'b0110;
assign label[15] = 4'b0100;
assign label[16] = 4'b0000;
assign label[17] = 4'b0100;
assign label[18] = 4'b0100;
assign label[19] = 4'b0011;
assign label[20] = 4'b0011;
assign label[21] = 4'b0001;
assign label[22] = 4'b0010;
assign label[23] = 4'b0111;
assign label[24] = 4'b0011;
assign label[25] = 4'b0100;
assign label[26] = 4'b1000;
assign label[27] = 4'b0101;
assign label[28] = 4'b1001;
assign label[29] = 4'b1000;
assign label[30] = 4'b0111;
assign label[31] = 4'b0110;
assign label[32] = 4'b0001;
assign label[33] = 4'b0001;
assign label[34] = 4'b0010;
assign label[35] = 4'b1000;
assign label[36] = 4'b0000;
assign label[37] = 4'b0111;
assign label[38] = 4'b0110;
assign label[39] = 4'b1001;
assign label[40] = 4'b0111;
assign label[41] = 4'b0011;
assign label[42] = 4'b0001;
assign label[43] = 4'b0000;
assign label[44] = 4'b1001;
assign label[45] = 4'b0011;
assign label[46] = 4'b0100;
assign label[47] = 4'b0010;
assign label[48] = 4'b0010;
assign label[49] = 4'b1000;
assign label[50] = 4'b0010;
assign label[51] = 4'b0111;
assign label[52] = 4'b0110;
assign label[53] = 4'b0100;
assign label[54] = 4'b0000;
assign label[55] = 4'b0100;
assign label[56] = 4'b0011;
assign label[57] = 4'b1001;
assign label[58] = 4'b0010;
assign label[59] = 4'b1000;
assign label[60] = 4'b0001;
assign label[61] = 4'b0011;
assign label[62] = 4'b0001;
assign label[63] = 4'b0011;
assign label[64] = 4'b0100;
assign label[65] = 4'b1001;
assign label[66] = 4'b0110;
assign label[67] = 4'b0100;
assign label[68] = 4'b0001;
assign label[69] = 4'b0100;
assign label[70] = 4'b0101;
assign label[71] = 4'b0101;
assign label[72] = 4'b0001;
assign label[73] = 4'b0011;
assign label[74] = 4'b1000;
assign label[75] = 4'b0001;
assign label[76] = 4'b0100;
assign label[77] = 4'b1000;
assign label[78] = 4'b1000;
assign label[79] = 4'b0001;
assign label[80] = 4'b0000;
assign label[81] = 4'b0101;
assign label[82] = 4'b0001;
assign label[83] = 4'b1001;
assign label[84] = 4'b0001;
assign label[85] = 4'b0010;
assign label[86] = 4'b0000;
assign label[87] = 4'b0100;
assign label[88] = 4'b0100;
assign label[89] = 4'b0110;
assign label[90] = 4'b0111;
assign label[91] = 4'b0111;
assign label[92] = 4'b0001;
assign label[93] = 4'b0111;
assign label[94] = 4'b1000;
assign label[95] = 4'b1000;
assign label[96] = 4'b0001;
assign label[97] = 4'b0010;
assign label[98] = 4'b0101;
assign label[99] = 4'b0001;
assign label[100] = 4'b1001;
assign label[101] = 4'b0000;
assign label[102] = 4'b0110;
assign label[103] = 4'b1001;
assign label[104] = 4'b0100;
assign label[105] = 4'b0111;
assign label[106] = 4'b0011;
assign label[107] = 4'b0001;
assign label[108] = 4'b0101;
assign label[109] = 4'b0101;
assign label[110] = 4'b1000;
assign label[111] = 4'b0010;
assign label[112] = 4'b0000;
assign label[113] = 4'b1001;
assign label[114] = 4'b0001;
assign label[115] = 4'b0011;
assign label[116] = 4'b0000;
assign label[117] = 4'b0110;
assign label[118] = 4'b0011;
assign label[119] = 4'b1000;
assign label[120] = 4'b0111;
assign label[121] = 4'b0000;
assign label[122] = 4'b0001;
assign label[123] = 4'b0110;
assign label[124] = 4'b0001;
assign label[125] = 4'b0010;
assign label[126] = 4'b0011;
assign label[127] = 4'b0110;
assign label[128] = 4'b0110;
assign label[129] = 4'b0111;
assign label[130] = 4'b0001;
assign label[131] = 4'b1001;
assign label[132] = 4'b0000;
assign label[133] = 4'b0100;
assign label[134] = 4'b0110;
assign label[135] = 4'b0010;
assign label[136] = 4'b0010;
assign label[137] = 4'b0111;
assign label[138] = 4'b0010;
assign label[139] = 4'b1001;
assign label[140] = 4'b0000;
assign label[141] = 4'b0000;
assign label[142] = 4'b1001;
assign label[143] = 4'b0010;
assign label[144] = 4'b0010;
assign label[145] = 4'b0001;
assign label[146] = 4'b0101;
assign label[147] = 4'b0110;
assign label[148] = 4'b1001;
assign label[149] = 4'b0110;
assign label[150] = 4'b0010;
assign label[151] = 4'b0011;
assign label[152] = 4'b0011;
assign label[153] = 4'b0111;
assign label[154] = 4'b1000;
assign label[155] = 4'b0100;
assign label[156] = 4'b0001;
assign label[157] = 4'b0010;
assign label[158] = 4'b0110;
assign label[159] = 4'b0110;
assign label[160] = 4'b0001;
assign label[161] = 4'b0010;
assign label[162] = 4'b1001;
assign label[163] = 4'b0111;
assign label[164] = 4'b1000;
assign label[165] = 4'b0101;
assign label[166] = 4'b0110;
assign label[167] = 4'b0001;
assign label[168] = 4'b0000;
assign label[169] = 4'b0011;
assign label[170] = 4'b0111;
assign label[171] = 4'b1001;
assign label[172] = 4'b0001;
assign label[173] = 4'b0011;
assign label[174] = 4'b0101;
assign label[175] = 4'b0010;
assign label[176] = 4'b0111;
assign label[177] = 4'b0101;
assign label[178] = 4'b0000;
assign label[179] = 4'b0001;
assign label[180] = 4'b0010;
assign label[181] = 4'b0010;
assign label[182] = 4'b0100;
assign label[183] = 4'b0111;
assign label[184] = 4'b0110;
assign label[185] = 4'b0111;
assign label[186] = 4'b1000;
assign label[187] = 4'b0110;
assign label[188] = 4'b0010;
assign label[189] = 4'b0011;
assign label[190] = 4'b1001;
assign label[191] = 4'b1000;
assign label[192] = 4'b0001;
assign label[193] = 4'b1001;
assign label[194] = 4'b0101;
assign label[195] = 4'b1000;
assign label[196] = 4'b0001;
assign label[197] = 4'b0001;
assign label[198] = 4'b0111;
assign label[199] = 4'b0010;
assign label[200] = 4'b1000;
assign label[201] = 4'b0110;
assign label[202] = 4'b1000;
assign label[203] = 4'b1000;
assign label[204] = 4'b1000;
assign label[205] = 4'b0011;
assign label[206] = 4'b0001;
assign label[207] = 4'b0111;
assign label[208] = 4'b0011;
assign label[209] = 4'b1000;
assign label[210] = 4'b0111;
assign label[211] = 4'b0000;
assign label[212] = 4'b0011;
assign label[213] = 4'b1001;
assign label[214] = 4'b0001;
assign label[215] = 4'b0110;
assign label[216] = 4'b0100;
assign label[217] = 4'b1000;
assign label[218] = 4'b0100;
assign label[219] = 4'b0010;
assign label[220] = 4'b0000;
assign label[221] = 4'b1001;
assign label[222] = 4'b0011;
assign label[223] = 4'b0011;
assign label[224] = 4'b0101;
assign label[225] = 4'b0101;
assign label[226] = 4'b1000;
assign label[227] = 4'b0110;
assign label[228] = 4'b0010;
assign label[229] = 4'b0011;
assign label[230] = 4'b1001;
assign label[231] = 4'b0101;
assign label[232] = 4'b0111;
assign label[233] = 4'b0101;
assign label[234] = 4'b1000;
assign label[235] = 4'b0111;
assign label[236] = 4'b0101;
assign label[237] = 4'b0001;
assign label[238] = 4'b0000;
assign label[239] = 4'b0100;
assign label[240] = 4'b0000;
assign label[241] = 4'b0010;
assign label[242] = 4'b0110;
assign label[243] = 4'b0111;
assign label[244] = 4'b1000;
assign label[245] = 4'b0101;
assign label[246] = 4'b1001;
assign label[247] = 4'b0100;
assign label[248] = 4'b0010;
assign label[249] = 4'b0001;
assign label[250] = 4'b1000;
assign label[251] = 4'b0100;
assign label[252] = 4'b1000;
assign label[253] = 4'b0011;
assign label[254] = 4'b0110;
assign label[255] = 4'b0010;
assign label[256] = 4'b1001;
assign label[257] = 4'b0110;
assign label[258] = 4'b1000;
assign label[259] = 4'b0001;
assign label[260] = 4'b0111;
assign label[261] = 4'b0000;
assign label[262] = 4'b0111;
assign label[263] = 4'b1001;
assign label[264] = 4'b0101;
assign label[265] = 4'b0110;
assign label[266] = 4'b0110;
assign label[267] = 4'b0000;
assign label[268] = 4'b0001;
assign label[269] = 4'b0000;
assign label[270] = 4'b0101;
assign label[271] = 4'b0110;
assign label[272] = 4'b0000;
assign label[273] = 4'b0111;
assign label[274] = 4'b0111;
assign label[275] = 4'b0111;
assign label[276] = 4'b1000;
assign label[277] = 4'b0011;
assign label[278] = 4'b0111;
assign label[279] = 4'b0001;
assign label[280] = 4'b0001;
assign label[281] = 4'b0011;
assign label[282] = 4'b0101;
assign label[283] = 4'b0001;
assign label[284] = 4'b1000;
assign label[285] = 4'b0100;
assign label[286] = 4'b0110;
assign label[287] = 4'b0100;
assign label[288] = 4'b1001;
assign label[289] = 4'b0001;
assign label[290] = 4'b0111;
assign label[291] = 4'b0101;
assign label[292] = 4'b0101;
assign label[293] = 4'b0011;
assign label[294] = 4'b0111;
assign label[295] = 4'b0010;
assign label[296] = 4'b1001;
assign label[297] = 4'b0110;
assign label[298] = 4'b0100;
assign label[299] = 4'b0101;
assign label[300] = 4'b1001;
assign label[301] = 4'b0110;
assign label[302] = 4'b0011;
assign label[303] = 4'b0011;
assign label[304] = 4'b1000;
assign label[305] = 4'b0110;
assign label[306] = 4'b0110;
assign label[307] = 4'b0111;
assign label[308] = 4'b0010;
assign label[309] = 4'b0010;
assign label[310] = 4'b0000;
assign label[311] = 4'b0001;
assign label[312] = 4'b0011;
assign label[313] = 4'b0011;
assign label[314] = 4'b0001;
assign label[315] = 4'b0111;
assign label[316] = 4'b1001;
assign label[317] = 4'b0000;
assign label[318] = 4'b0010;
assign label[319] = 4'b0101;
assign label[320] = 4'b0110;
assign label[321] = 4'b0001;
assign label[322] = 4'b0111;
assign label[323] = 4'b1000;
assign label[324] = 4'b0001;
assign label[325] = 4'b0001;
assign label[326] = 4'b0110;
assign label[327] = 4'b1000;
assign label[328] = 4'b0000;
assign label[329] = 4'b0000;
assign label[330] = 4'b0101;
assign label[331] = 4'b0001;
assign label[332] = 4'b0010;
assign label[333] = 4'b0111;
assign label[334] = 4'b0110;
assign label[335] = 4'b0010;
assign label[336] = 4'b0100;
assign label[337] = 4'b1001;
assign label[338] = 4'b1001;
assign label[339] = 4'b0001;
assign label[340] = 4'b0100;
assign label[341] = 4'b0101;
assign label[342] = 4'b0001;
assign label[343] = 4'b1000;
assign label[344] = 4'b0010;
assign label[345] = 4'b0110;
assign label[346] = 4'b0111;
assign label[347] = 4'b1001;
assign label[348] = 4'b0010;
assign label[349] = 4'b0100;
assign label[350] = 4'b0110;
assign label[351] = 4'b0111;
assign label[352] = 4'b0011;
assign label[353] = 4'b0110;
assign label[354] = 4'b0101;
assign label[355] = 4'b0101;
assign label[356] = 4'b1001;
assign label[357] = 4'b0010;
assign label[358] = 4'b0101;
assign label[359] = 4'b0111;
assign label[360] = 4'b0010;
assign label[361] = 4'b0001;
assign label[362] = 4'b0011;
assign label[363] = 4'b0011;
assign label[364] = 4'b0110;
assign label[365] = 4'b1000;
assign label[366] = 4'b0101;
assign label[367] = 4'b0000;
assign label[368] = 4'b1001;
assign label[369] = 4'b0001;
assign label[370] = 4'b0000;
assign label[371] = 4'b0011;
assign label[372] = 4'b0101;
assign label[373] = 4'b0010;
assign label[374] = 4'b0101;
assign label[375] = 4'b0110;
assign label[376] = 4'b0000;
assign label[377] = 4'b0010;
assign label[378] = 4'b0001;
assign label[379] = 4'b0001;
assign label[380] = 4'b0111;
assign label[381] = 4'b0000;
assign label[382] = 4'b0000;
assign label[383] = 4'b0000;
assign label[384] = 4'b0000;
assign label[385] = 4'b0001;
assign label[386] = 4'b0011;
assign label[387] = 4'b0110;
assign label[388] = 4'b0010;
assign label[389] = 4'b0110;
assign label[390] = 4'b1001;
assign label[391] = 4'b0101;
assign label[392] = 4'b1001;
assign label[393] = 4'b0101;
assign label[394] = 4'b0100;
assign label[395] = 4'b0000;
assign label[396] = 4'b0001;
assign label[397] = 4'b0110;
assign label[398] = 4'b0110;
assign label[399] = 4'b0110;
assign label[400] = 4'b1000;
assign label[401] = 4'b1000;
assign label[402] = 4'b1000;
assign label[403] = 4'b0001;
assign label[404] = 4'b1000;
assign label[405] = 4'b1000;
assign label[406] = 4'b1001;
assign label[407] = 4'b0100;
assign label[408] = 4'b0001;
assign label[409] = 4'b0111;
assign label[410] = 4'b1000;
assign label[411] = 4'b1000;
assign label[412] = 4'b0001;
assign label[413] = 4'b0000;
assign label[414] = 4'b0000;
assign label[415] = 4'b0110;
assign label[416] = 4'b0011;
assign label[417] = 4'b0100;
assign label[418] = 4'b0000;
assign label[419] = 4'b0001;
assign label[420] = 4'b0111;
assign label[421] = 4'b0101;
assign label[422] = 4'b0110;
assign label[423] = 4'b0001;
assign label[424] = 4'b0001;
assign label[425] = 4'b0111;
assign label[426] = 4'b0100;
assign label[427] = 4'b0110;
assign label[428] = 4'b0001;
assign label[429] = 4'b0010;
assign label[430] = 4'b1001;
assign label[431] = 4'b1000;
assign label[432] = 4'b0110;
assign label[433] = 4'b0010;
assign label[434] = 4'b1000;
assign label[435] = 4'b1000;
assign label[436] = 4'b0001;
assign label[437] = 4'b0001;
assign label[438] = 4'b0001;
assign label[439] = 4'b0011;
assign label[440] = 4'b1000;
assign label[441] = 4'b0101;
assign label[442] = 4'b0101;
assign label[443] = 4'b1000;
assign label[444] = 4'b0000;
assign label[445] = 4'b0101;
assign label[446] = 4'b1001;
assign label[447] = 4'b0000;
assign label[448] = 4'b0010;
assign label[449] = 4'b0000;
assign label[450] = 4'b0111;
assign label[451] = 4'b0101;
assign label[452] = 4'b1000;
assign label[453] = 4'b0011;
assign label[454] = 4'b0000;
assign label[455] = 4'b0010;
assign label[456] = 4'b1000;
assign label[457] = 4'b0110;
assign label[458] = 4'b0110;
assign label[459] = 4'b0011;
assign label[460] = 4'b0000;
assign label[461] = 4'b0100;
assign label[462] = 4'b0100;
assign label[463] = 4'b0110;
assign label[464] = 4'b0110;
assign label[465] = 4'b1000;
assign label[466] = 4'b0110;
assign label[467] = 4'b0001;
assign label[468] = 4'b0110;
assign label[469] = 4'b0000;
assign label[470] = 4'b0111;
assign label[471] = 4'b0100;
assign label[472] = 4'b1001;
assign label[473] = 4'b0111;
assign label[474] = 4'b1000;
assign label[475] = 4'b1001;
assign label[476] = 4'b0010;
assign label[477] = 4'b1001;
assign label[478] = 4'b0111;
assign label[479] = 4'b0000;
assign label[480] = 4'b0011;
assign label[481] = 4'b0111;
assign label[482] = 4'b1000;
assign label[483] = 4'b0111;
assign label[484] = 4'b0111;
assign label[485] = 4'b0111;
assign label[486] = 4'b1000;
assign label[487] = 4'b0011;
assign label[488] = 4'b0111;
assign label[489] = 4'b0011;
assign label[490] = 4'b0001;
assign label[491] = 4'b0001;
assign label[492] = 4'b0110;
assign label[493] = 4'b0010;
assign label[494] = 4'b0111;
assign label[495] = 4'b0110;
assign label[496] = 4'b1000;
assign label[497] = 4'b0000;
assign label[498] = 4'b0110;
assign label[499] = 4'b0010;
assign label[500] = 4'b0000;
assign label[501] = 4'b1000;
assign label[502] = 4'b1000;
assign label[503] = 4'b0111;
assign label[504] = 4'b1001;
assign label[505] = 4'b1001;
assign label[506] = 4'b1000;
assign label[507] = 4'b0101;
assign label[508] = 4'b0101;
assign label[509] = 4'b0100;
assign label[510] = 4'b0100;
assign label[511] = 4'b0110;
assign label[512] = 4'b0011;
assign label[513] = 4'b0111;
assign label[514] = 4'b0110;
assign label[515] = 4'b1000;
assign label[516] = 4'b0001;
assign label[517] = 4'b0011;
assign label[518] = 4'b0111;
assign label[519] = 4'b0100;
assign label[520] = 4'b0010;
assign label[521] = 4'b0011;
assign label[522] = 4'b0001;
assign label[523] = 4'b0101;
assign label[524] = 4'b0011;
assign label[525] = 4'b1000;
assign label[526] = 4'b0001;
assign label[527] = 4'b0110;
assign label[528] = 4'b0101;
assign label[529] = 4'b0100;
assign label[530] = 4'b0001;
assign label[531] = 4'b0000;
assign label[532] = 4'b0010;
assign label[533] = 4'b0111;
assign label[534] = 4'b1000;
assign label[535] = 4'b0011;
assign label[536] = 4'b0110;
assign label[537] = 4'b0111;
assign label[538] = 4'b0111;
assign label[539] = 4'b0011;
assign label[540] = 4'b0001;
assign label[541] = 4'b0100;
assign label[542] = 4'b0101;
assign label[543] = 4'b0010;
assign label[544] = 4'b0011;
assign label[545] = 4'b0001;
assign label[546] = 4'b0111;
assign label[547] = 4'b0010;
assign label[548] = 4'b1001;
assign label[549] = 4'b0001;
assign label[550] = 4'b0100;
assign label[551] = 4'b0111;
assign label[552] = 4'b0010;
assign label[553] = 4'b1001;
assign label[554] = 4'b1001;
assign label[555] = 4'b0010;
assign label[556] = 4'b0011;
assign label[557] = 4'b0111;
assign label[558] = 4'b0010;
assign label[559] = 4'b0110;
assign label[560] = 4'b0011;
assign label[561] = 4'b0000;
assign label[562] = 4'b0001;
assign label[563] = 4'b0111;
assign label[564] = 4'b0010;
assign label[565] = 4'b1001;
assign label[566] = 4'b1001;
assign label[567] = 4'b0011;
assign label[568] = 4'b0011;
assign label[569] = 4'b0000;
assign label[570] = 4'b0101;
assign label[571] = 4'b0111;
assign label[572] = 4'b0000;
assign label[573] = 4'b0011;
assign label[574] = 4'b0011;
assign label[575] = 4'b0110;
assign label[576] = 4'b0010;
assign label[577] = 4'b0111;
assign label[578] = 4'b0110;
assign label[579] = 4'b0011;
assign label[580] = 4'b0100;
assign label[581] = 4'b0001;
assign label[582] = 4'b0001;
assign label[583] = 4'b0101;
assign label[584] = 4'b0000;
assign label[585] = 4'b0100;
assign label[586] = 4'b0110;
assign label[587] = 4'b1000;
assign label[588] = 4'b0110;
assign label[589] = 4'b0100;
assign label[590] = 4'b0100;
assign label[591] = 4'b0100;
assign label[592] = 4'b0011;
assign label[593] = 4'b0110;
assign label[594] = 4'b0000;
assign label[595] = 4'b0110;
assign label[596] = 4'b0001;
assign label[597] = 4'b0111;
assign label[598] = 4'b0111;
assign label[599] = 4'b0110;
assign label[600] = 4'b0100;
assign label[601] = 4'b0011;
assign label[602] = 4'b0000;
assign label[603] = 4'b0011;
assign label[604] = 4'b0000;
assign label[605] = 4'b0101;
assign label[606] = 4'b0010;
assign label[607] = 4'b0100;
assign label[608] = 4'b0111;
assign label[609] = 4'b0110;
assign label[610] = 4'b0011;
assign label[611] = 4'b0000;
assign label[612] = 4'b1000;
assign label[613] = 4'b0110;
assign label[614] = 4'b0111;
assign label[615] = 4'b0001;
assign label[616] = 4'b0100;
assign label[617] = 4'b0100;
assign label[618] = 4'b0011;
assign label[619] = 4'b0101;
assign label[620] = 4'b1000;
assign label[621] = 4'b0010;
assign label[622] = 4'b0110;
assign label[623] = 4'b1000;
assign label[624] = 4'b0011;
assign label[625] = 4'b0111;
assign label[626] = 4'b1001;
assign label[627] = 4'b0000;
assign label[628] = 4'b0010;
assign label[629] = 4'b0000;
assign label[630] = 4'b0110;
assign label[631] = 4'b0000;
assign label[632] = 4'b0110;
assign label[633] = 4'b1000;
assign label[634] = 4'b0111;
assign label[635] = 4'b0100;
assign label[636] = 4'b0010;
assign label[637] = 4'b0101;
assign label[638] = 4'b1001;
assign label[639] = 4'b0000;
assign label[640] = 4'b0011;
assign label[641] = 4'b0011;
assign label[642] = 4'b1001;
assign label[643] = 4'b0001;
assign label[644] = 4'b0011;
assign label[645] = 4'b0110;
assign label[646] = 4'b0000;
assign label[647] = 4'b0110;
assign label[648] = 4'b0001;
assign label[649] = 4'b0101;
assign label[650] = 4'b1000;
assign label[651] = 4'b0100;
assign label[652] = 4'b0010;
assign label[653] = 4'b1001;
assign label[654] = 4'b0001;
assign label[655] = 4'b0111;
assign label[656] = 4'b1001;
assign label[657] = 4'b0110;
assign label[658] = 4'b1001;
assign label[659] = 4'b0001;
assign label[660] = 4'b0000;
assign label[661] = 4'b0110;
assign label[662] = 4'b0101;
assign label[663] = 4'b0100;
assign label[664] = 4'b0011;
assign label[665] = 4'b1001;
assign label[666] = 4'b0111;
assign label[667] = 4'b0010;
assign label[668] = 4'b0110;
assign label[669] = 4'b0011;
assign label[670] = 4'b0110;
assign label[671] = 4'b0111;
assign label[672] = 4'b0010;
assign label[673] = 4'b0011;
assign label[674] = 4'b0000;
assign label[675] = 4'b0000;
assign label[676] = 4'b0010;
assign label[677] = 4'b0000;
assign label[678] = 4'b0101;
assign label[679] = 4'b1001;
assign label[680] = 4'b0111;
assign label[681] = 4'b0100;
assign label[682] = 4'b0101;
assign label[683] = 4'b0000;
assign label[684] = 4'b0001;
assign label[685] = 4'b0111;
assign label[686] = 4'b0110;
assign label[687] = 4'b0010;
assign label[688] = 4'b1000;
assign label[689] = 4'b0110;
assign label[690] = 4'b1000;
assign label[691] = 4'b1000;
assign label[692] = 4'b0110;
assign label[693] = 4'b1001;
assign label[694] = 4'b0010;
assign label[695] = 4'b0110;
assign label[696] = 4'b0000;
assign label[697] = 4'b0000;
assign label[698] = 4'b1000;
assign label[699] = 4'b0000;
assign label[700] = 4'b0000;
assign label[701] = 4'b0111;
assign label[702] = 4'b1001;
assign label[703] = 4'b0111;
assign label[704] = 4'b0100;
assign label[705] = 4'b1000;
assign label[706] = 4'b1001;
assign label[707] = 4'b1001;
assign label[708] = 4'b1000;
assign label[709] = 4'b0101;
assign label[710] = 4'b1000;
assign label[711] = 4'b1001;
assign label[712] = 4'b0000;
assign label[713] = 4'b0010;
assign label[714] = 4'b1001;
assign label[715] = 4'b0110;
assign label[716] = 4'b0111;
assign label[717] = 4'b1000;
assign label[718] = 4'b0110;
assign label[719] = 4'b0101;
assign label[720] = 4'b0110;
assign label[721] = 4'b0011;
assign label[722] = 4'b0101;
assign label[723] = 4'b0010;
assign label[724] = 4'b0010;
assign label[725] = 4'b0010;
assign label[726] = 4'b1000;
assign label[727] = 4'b0111;
assign label[728] = 4'b0010;
assign label[729] = 4'b0101;
assign label[730] = 4'b0110;
assign label[731] = 4'b0010;
assign label[732] = 4'b0011;
assign label[733] = 4'b0001;
assign label[734] = 4'b0010;
assign label[735] = 4'b1001;
assign label[736] = 4'b0110;
assign label[737] = 4'b0011;
assign label[738] = 4'b0001;
assign label[739] = 4'b0011;
assign label[740] = 4'b0000;
assign label[741] = 4'b0101;
assign label[742] = 4'b1000;
assign label[743] = 4'b0001;
assign label[744] = 4'b0110;
assign label[745] = 4'b1001;
assign label[746] = 4'b0000;
assign label[747] = 4'b0011;
assign label[748] = 4'b0000;
assign label[749] = 4'b0001;

    always @(*)
    begin
        if (read_input == 1'b1)
            out = label[addr];
        else
            out = 4'bZ;
    end

endmodule   


`timescale 1ns/1ns
module camparator(input[3:0] in1, in2, output eq);

assign eq = (in1 == in2); 

endmodule
